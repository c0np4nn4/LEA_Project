module LEA_BlockSubtractor_tb;

reg [31:0] A;
reg [31:0] B;
wire [31:0] Result;

LEA_BlockSubtractor
 U0 (
  .A(A),
  .B(B),
  .Result(Result));

  initial
  begin
    A = 32'b10100011111100110111101011111000;
    #100 A = 32'b01101010101001110011100100011010;
    #100 A = 32'b00100110110111111100001101011110;
    #100 A = 32'b01101010110110110010101111011010;
    #100 A = 32'b11111101101101111111110100100000;
    #100 A = 32'b10110000110100111110011100010001;
    #100 A = 32'b11110010001011000111110111011111;
    #100 A = 32'b10101101011100110000100010100111;
    #100 A = 32'b11011010101110000100001001111000;
    #100 A = 32'b00001011001110111110011000110110;
    #100 A = 32'b11011011000010110001110010011010;
    #100 A = 32'b11010110011110111100000001110111;
    #100 A = 32'b00111010010000001110011101010011;
    #100 A = 32'b11110010100101000111010010011110;
    #100 A = 32'b00000101010010100111000001110111;
    #100 A = 32'b01011011000000000100010000111110;
    #100 A = 32'b01110010001111111001101000101100;
    #100 A = 32'b00001110000001101111010001100111;
    #100 A = 32'b10010001000100110101010001101011;
    #100 A = 32'b11100010110000001110101100010110;
    #100 A = 32'b01011010011011100100110110100010;
    #100 A = 32'b10100001001000111101111000101010;
    #100 A = 32'b10000011100100101000010111010001;
    #100 A = 32'b10001010110100100110110010100111;
    #100 A = 32'b00011101001111010110010111010111;
    #100 A = 32'b11010100010001000001011001010011;
    #100 A = 32'b10010001001001110111010111111110;
    #100 A = 32'b10101001000000011010001000110010;
    #100 A = 32'b11110001110000111111000110100000;
    #100 A = 32'b11101011101010100010000000111011;
    #100 A = 32'b01101001010100000110110111111111;
    #100 A = 32'b11001111111111100001010101011010;
    #100 A = 32'b01001010011000100101110000110001;
    #100 A = 32'b00110011011100101010110010000001;
    #100 A = 32'b01110011011001111110000001010101;
    #100 A = 32'b01011000010100110110110111001010;
    #100 A = 32'b00010001110111101110011001110001;
    #100 A = 32'b10000011000100011111000100110111;
    #100 A = 32'b11010000001101111110101000100101;
    #100 A = 32'b11110101011000100011010010101011;
    #100 A = 32'b11111001111100110001010000010000;
    #100 A = 32'b11110010000001101000100000000010;
    #100 A = 32'b00000100100101010000010111110100;
    #100 A = 32'b10000000010010100001010000101110;
    #100 A = 32'b10110111111001111010001000100000;
    #100 A = 32'b11111110101101011001001111101000;
    #100 A = 32'b10110000000100011001111011110110;
    #100 A = 32'b10011110001001111001010001011000;
    #100 A = 32'b11100001001011010000001010101101;
    #100 A = 32'b10000100001101010010011101110000;
    #100 A = 32'b01111010000110111100101010000111;
    #100 A = 32'b00100001011111000011111011110110;
    #100 A = 32'b11011001110111100011111110101100;
    #100 A = 32'b00111000111000110101101101011110;
    #100 A = 32'b00000110011101000001010010000100;
    #100 A = 32'b00001010001011011000101110111101;
    #100 A = 32'b01010000000011100001111101100001;
    #100 A = 32'b01111010110110110011011001000000;
    #100 A = 32'b00010010100100110101100110011011;
    #100 A = 32'b01100010011110101011011010010110;
    #100 A = 32'b01100001111110001001101101100111;
    #100 A = 32'b10100001110100101010101101101111;
    #100 A = 32'b01110001010001101101100001111111;
    #100 A = 32'b10000011000100001010111011111111;
    #100 A = 32'b01111111100011001100000010101111;
    #100 A = 32'b00010000110111010100010011101110;
    #100 A = 32'b10011001110101011111010110100110;
    #100 A = 32'b11101101100110100000000010000110;
    #100 A = 32'b11000011011011001100011100010010;
    #100 A = 32'b11111101010100011110101111111100;
    #100 A = 32'b01101010001000100000000000111010;
    #100 A = 32'b11101011001010110100001010111010;
    #100 A = 32'b00010100010010100101001000001111;
    #100 A = 32'b11011001010010001010100101001110;
    #100 A = 32'b11101000011001011011010111100110;
    #100 A = 32'b10001110111001101000111111100111;
    #100 A = 32'b11111000100011101111101111111101;
    #100 A = 32'b00100000011110100000111000000000;
    #100 A = 32'b00100010101111011000011011101011;
    #100 A = 32'b01000110111100001110001001011011;
    #100 A = 32'b10100111111101010011100011000010;
    #100 A = 32'b00000011110111001011010101111001;
    #100 A = 32'b11110011010001000001110001100101;
    #100 A = 32'b10000000100000010001010101111100;
    #100 A = 32'b00101011110110111110110100000010;
    #100 A = 32'b11101101100101001101001011010010;
    #100 A = 32'b11110111000110000101001011010111;
    #100 A = 32'b01110111010000100000001111011111;
    #100 A = 32'b01100100100010100000011100011000;
    #100 A = 32'b11101100000001101111101111100000;
    #100 A = 32'b00110001101101011001000100111111;
    #100 A = 32'b10011011000110000001101110110101;
    #100 A = 32'b10110000110100001101101110011000;
    #100 A = 32'b01100101110000000000001101010111;
    #100 A = 32'b00101111011110101011001110000010;
    #100 A = 32'b10100000010111101011110100100001;
    #100 A = 32'b01100011101011010100110100111000;
    #100 A = 32'b01100000010010101010110101111111;
    #100 A = 32'b11101100001111000000010110001101;
    #100 A = 32'b11100110111000101100100110111010;
  end

  initial
  begin
    B = 32'b01011011111101110101110111110011;
    #100 B = 32'b00000111111110011000000001001101;
    #100 B = 32'b00111110001000111110010010111010;
    #100 B = 32'b00011111111000100110010100001010;
    #100 B = 32'b01001011111000010100001101111011;
    #100 B = 32'b00100100101000101100011101000001;
    #100 B = 32'b10010011011010011011000011010011;
    #100 B = 32'b01011111010000100001011100111011;
    #100 B = 32'b10011101101100001001101111011001;
    #100 B = 32'b11100010101100001111111100000011;
    #100 B = 32'b10100001001010100001001011100100;
    #100 B = 32'b11110000001001011001100011110101;
    #100 B = 32'b00010001011100000000001100010000;
    #100 B = 32'b01111101001000101010000101111001;
    #100 B = 32'b10001101001110001110010010001001;
    #100 B = 32'b00111001110011101110100010110111;
    #100 B = 32'b11001110100110000001001001110010;
    #100 B = 32'b11001110100111011110010100001000;
    #100 B = 32'b10010100011000001100100011001010;
    #100 B = 32'b00010111011010001011010101110011;
    #100 B = 32'b00011000000011100110010110010000;
    #100 B = 32'b01000100111101001110101111010101;
    #100 B = 32'b00010101001100011100100101011111;
    #100 B = 32'b10001001011110110100111010001010;
    #100 B = 32'b01011010011001110010000011111000;
    #100 B = 32'b00111000000110010100010010101000;
    #100 B = 32'b11110111110011010100000000110011;
    #100 B = 32'b01100000001101001101101001100110;
    #100 B = 32'b01001111010100101101110010110011;
    #100 B = 32'b00001001101000001001001000011000;
    #100 B = 32'b10111000001011000110101110101001;
    #100 B = 32'b10101001001111100110111100101011;
    #100 B = 32'b11010101010010000111001100001011;
    #100 B = 32'b10111110100100011110100001111101;
    #100 B = 32'b00111110110000111111010101001101;
    #100 B = 32'b01111001100010111001011011011110;
    #100 B = 32'b10110110010110110100110001110011;
    #100 B = 32'b11000110100100100001001000110110;
    #100 B = 32'b01001111101110001111000010000000;
    #100 B = 32'b10101001011111001001001111100011;
    #100 B = 32'b11001100010110101100101001000010;
    #100 B = 32'b00001101011001000111111011000001;
    #100 B = 32'b01010000111010010101000001010100;
    #100 B = 32'b00101011111001101111001001111101;
    #100 B = 32'b01100110110110000111001111100001;
    #100 B = 32'b11111101001000001110000101000110;
    #100 B = 32'b11100111001110110100001100101000;
    #100 B = 32'b10001011101101111000001000100000;
    #100 B = 32'b10100110001001011011000100000011;
    #100 B = 32'b11110001100010100100010001011010;
    #100 B = 32'b01101000010111101111000111100100;
    #100 B = 32'b01010010110010111110001001100001;
    #100 B = 32'b01110100100100111110011100011111;
    #100 B = 32'b11011010111101111101100001101111;
    #100 B = 32'b10001001001000100011000110001101;
    #100 B = 32'b01110000101001101110111001101001;
    #100 B = 32'b11011010111010101100010110110000;
    #100 B = 32'b11111010000100111111110010010010;
    #100 B = 32'b10010111101111011101010001001000;
    #100 B = 32'b01101010001001001100111101000010;
    #100 B = 32'b00010010000011110111010000000011;
    #100 B = 32'b00111001010011110110110110110011;
    #100 B = 32'b11101010100111110100111100100111;
    #100 B = 32'b00100001100100100100111001110110;
    #100 B = 32'b11111111111010110001111000110100;
    #100 B = 32'b01000100101101000000101011101000;
    #100 B = 32'b11000100101001001111110101101000;
    #100 B = 32'b10001100101101111001011010000001;
    #100 B = 32'b10111101110111011101001101011001;
    #100 B = 32'b11100010001111101001010100110101;
    #100 B = 32'b11011110101010010111110100010100;
    #100 B = 32'b01010101011010110010101011111001;
    #100 B = 32'b11000000011000000010010101001110;
    #100 B = 32'b00011101011100010111110001011110;
    #100 B = 32'b01101000010111110001110000111000;
    #100 B = 32'b10001001011000001100011011000000;
    #100 B = 32'b10100100110101100100110110001001;
    #100 B = 32'b01101000110000010110010100011110;
    #100 B = 32'b11000111110010101100101010100111;
    #100 B = 32'b00110110111010010010100100101111;
    #100 B = 32'b00100010001111000110100110110110;
    #100 B = 32'b01111001010011011111000011111011;
    #100 B = 32'b10101111010111101111101110101100;
    #100 B = 32'b00001001110101000110100101000010;
    #100 B = 32'b11010010101001110101010010011110;
    #100 B = 32'b00100101010000011001001101000000;
    #100 B = 32'b11111000010001011101001101101110;
    #100 B = 32'b11111110111011011110011110111011;
    #100 B = 32'b01000000100111010001111110010101;
    #100 B = 32'b11001111101011010001100000110001;
    #100 B = 32'b11101000011101101101000110110100;
    #100 B = 32'b00000001001111111001010011010010;
    #100 B = 32'b11100110110100000011000010010111;
    #100 B = 32'b11100100111101101101010010101110;
    #100 B = 32'b00000011101010111100000100100011;
    #100 B = 32'b01000011110101110101101001000101;
    #100 B = 32'b00100000001111110000000111011110;
    #100 B = 32'b00101011100011111011000000001011;
    #100 B = 32'b11100101011111001001110010011001;
    #100 B = 32'b01010101010011101111110111000000;
  end

endmodule
