module LEA_128BitsDivideIn16x8Register_tb;

reg [127:0] Din;
wire [7:0] Dout0;
wire [7:0] Dout1;
wire [7:0] Dout10;
wire [7:0] Dout11;
wire [7:0] Dout12;
wire [7:0] Dout13;
wire [7:0] Dout14;
wire [7:0] Dout15;
wire [7:0] Dout2;
wire [7:0] Dout3;
wire [7:0] Dout4;
wire [7:0] Dout5;
wire [7:0] Dout6;
wire [7:0] Dout7;
wire [7:0] Dout8;
wire [7:0] Dout9;

LEA_128BitsDivideIn16x8Register
 U0 (
  .Din(Din),
  .Dout0(Dout0),
  .Dout1(Dout1),
  .Dout10(Dout10),
  .Dout11(Dout11),
  .Dout12(Dout12),
  .Dout13(Dout13),
  .Dout14(Dout14),
  .Dout15(Dout15),
  .Dout2(Dout2),
  .Dout3(Dout3),
  .Dout4(Dout4),
  .Dout5(Dout5),
  .Dout6(Dout6),
  .Dout7(Dout7),
  .Dout8(Dout8),
  .Dout9(Dout9));

  initial
  begin
    Din = 128'b00111111011101110101100100101000111100110001001100111110110110110000110100111101101100011101010100001111001010011110100100101000;
    #100 Din = 128'b11111111111011001001101111101010000010000011010000000001010100000010001010111110110110000000110001100110101000001111110001100010;
    #100 Din = 128'b01100010011011010100110101011101010000111101111100000010101000110100100100000001101000101011011000101100111011011101101011011010;
    #100 Din = 128'b11100101100111000110011110011110101100000011110100111111111110110001000111010100111111011101001100011101100000010001101000001100;
    #100 Din = 128'b10110110000011010000000001111100101000011010001001010101000011111010001011011100111000000111111111011101100101110000011001111101;
    #100 Din = 128'b11111101000100100101110011001001101110011110110001000011110011010000011100011010111000001100001000001110001100010110100110010011;
    #100 Din = 128'b10000110010011110000111110001001000001110011101101000011001100011001100011110110110010011111010101011011111001100000111001010001;
    #100 Din = 128'b00010101000001010000011001000100100011001101101001000001001111000110010101110100010110110010100001001101100010110000100101011000;
    #100 Din = 128'b00011110100101010001010001010001101011111111100010101011010100100110101110101000011011001010011110100101010101001000000000111111;
    #100 Din = 128'b10010001101100010100111111011101110001010110101110110011001110110001101100011000011011100010101011100111110010011100001001001101;
    #100 Din = 128'b01111011111110011000110010101010011001000101100011011111101001001111011010001010100110100011101100110101111110001110011010110110;
    #100 Din = 128'b10010111010110110101101011011110010100011101110111010100100000101000010010110011101101011001011111111011011001110110110000000111;
    #100 Din = 128'b11111111100100000100100101111100010100000010000111111011100011101100100111011000100111010001011011011100110010110010000010010000;
    #100 Din = 128'b11111011101111100111110001010000100010011111100100111000111000010011011001000111100110001000011110100100101101101110111011100110;
    #100 Din = 128'b00111110010001111000010111011100101100000010110110100100001101011100001111001000001110000100100110000110001011111010011111100010;
    #100 Din = 128'b11110011000111001111000111100111001011111000011000110011011000011110100100000001010110100010101101010110101101010001110110000100;
    #100 Din = 128'b10110011101101000010111011101010111110101011011000011101001111101100001110011010101011111101011001011110111101010111000101000100;
    #100 Din = 128'b00101000111100110111000010001000101100000000101001111000010000010000111001101000100011111111010100110000010100110110101001101110;
    #100 Din = 128'b01000101110110000000101011111110110011100111011011010100110111100100100110101110110100110101010111101100111111000111110101110110;
    #100 Din = 128'b01011110011000001000111010100100100001010101100101011110101001010000000111000111001010010010010100011100111000011100001000100110;
    #100 Din = 128'b10110110100010111000010100001111010000110000000101001000001100110110101010010101111110110110101110000111100100000101000111001001;
    #100 Din = 128'b00100101110000011001000011011101111101110110111101011010010101101101010000001100011001110100011010101111101011001101111001110010;
    #100 Din = 128'b01010011010001000011111011010010111100011000011001001111111000010000010110111110110001011101000011011100111100000110010101011001;
    #100 Din = 128'b10000111011111101110011100111000001011110001110110001011111111101011010111000111001110111010001001010000111010101100101111001110;
    #100 Din = 128'b01111100001011000110001010100100110000100010001010111010110111010100110001010110001101101000101010011010101101101100011110001101;
    #100 Din = 128'b10011100001011001100001100000010101011000010110001011101111000011101101011001111110101011101111010011110111001100011001100110000;
    #100 Din = 128'b10000001111111101101001010010110010101111010001011101011110001010101011110100100110110111011111111111001010001010000110110111001;
    #100 Din = 128'b00100100011001100010000001111001110100101100110000110111010111100000000010010001101000111010100010100111011000111001001101101000;
    #100 Din = 128'b11110111001101010100101100010111010011001100110001010000111010000100111001111100011101000011110110111111011101000010001110110000;
    #100 Din = 128'b10100101101010100111000010101000101100100011100110011001000100010111111000101100000111010011101011101000111101110011100001010110;
    #100 Din = 128'b10111010010101011000101110011001101010001001101110100101000011111100111111101111001100010100001110101101110111011110010100101001;
    #100 Din = 128'b00100011111111010000011110000101111110110100101001000010101010011101111010001010010011100100111110111001110000011111010111000011;
    #100 Din = 128'b11100001010001100101110110111111100011000110001111001110100100110110101001000010001001111101101100010001011111010101101110110111;
    #100 Din = 128'b01011011111011011111001111000101000111110000011101010101101100001000000100010100111001110110000011100001011010100010011111000100;
    #100 Din = 128'b11010111100111111111001010000110011011010111010001100111110101010101010110000110100011101101100010000101100100111001101010111000;
    #100 Din = 128'b00010101110110000101100011000001101001100010110101100000000000010111001001011000001011110011100101001101110100000001001110001010;
    #100 Din = 128'b01010010011001001010011001111000000110101110010100111111011010010101100011011010000101001010000011001100100110111010100000110100;
    #100 Din = 128'b00111001000100010011111110111001000010111010010111001010000001110111100001001011000001010110111000011111010111011011011001110100;
    #100 Din = 128'b00101010001111101010000111001100100010101111100111011000110100010010011111100000101111110110101110100000101001101100001111010101;
    #100 Din = 128'b10001111000101000001011010001100111110110001010011111000010110100010011000010011111010111110010100011010001000100000011100011101;
    #100 Din = 128'b11100011001100010011111001000011111011101010010011110010001111100101011001110011110001001100001111011001011001100110101010110011;
    #100 Din = 128'b10110111001001010100100100111001010001011111100010010010101010101111001010010000110001001010111110011111011100110100100100011011;
    #100 Din = 128'b11011110010101010000110110100010000101111100000110001110111111100011110010110010110111001100001011101010001001000100111101110111;
    #100 Din = 128'b11100101110101101101100110101010111110000111111111000110100001100111101101100001010101011111010001011111110000100000011110000111;
    #100 Din = 128'b01100011111011001101000000010000000101110110011101010010110101010101001000010101011011011000001011000001110000111110111010111000;
    #100 Din = 128'b10000111001100111000111011111111110001111011000110001011110010100111000110001111100100000011111101010101000100000100110101110110;
    #100 Din = 128'b10011011110100011010101011010011010101111111111011000000110010100101101010000110111100110001110111100011010010111110111111110010;
    #100 Din = 128'b01110011010101110101011110100110001100010110100010001001001001101100001011101011111001011110100111010010101011010101111101110111;
    #100 Din = 128'b10000100000001011000101001011111110010001100101000100100010101101110111101010111111100110111101111001001001111011110001010011001;
    #100 Din = 128'b00011000100011001000111011101100001001111010111000111100110000001010110000101011001101101011110011110101110010110011101101101111;
    #100 Din = 128'b10111010101001110011110101001000001000100100010111110010101110111001100110011001111011110100000010101110001001101111000100010001;
    #100 Din = 128'b11100110100001001011010110111001110111111101110000000010110101100001100011011010011111011010100011011100010001100101010000110100;
    #100 Din = 128'b11010000001111101011011001101100001011110010011110011101011000101110001110010111110111011011010101111011101010001011101111100001;
    #100 Din = 128'b00011010011110001110111011101111000011001000000001101000111111111111101111010001010010101100101110010010000011101000110011001110;
    #100 Din = 128'b11011101001100101000111111111111001110101011100101001110001010100101011111100111100110010010100111000111111011001011010011100111;
    #100 Din = 128'b10100111010011111111001110110010001011111101001101010000101000111100100010110100000110001000001000000110010100110101001110100000;
    #100 Din = 128'b11100011000111101101111010101101111010111111011010110110100001100111100000101010000010000001111100110010010111100001110101010110;
    #100 Din = 128'b11000000000011101010001100010011110101010001001001110000011100010100000111101111111001111001000010000000110100100111110001010111;
    #100 Din = 128'b01011011011011100110011111101100000011101011011100111000111101101111011001001000011111110111001001101101010010011101000101011111;
    #100 Din = 128'b11001111011100010001111110001100010100011111000111111010001010111100011011001101011110001110100010111010110010001110110011011100;
    #100 Din = 128'b10010011011111110010111010110010011000010000101101101111100100001010110100110000110001000100111110011000111011001011100010011010;
    #100 Din = 128'b01100001100000101001010000100100000101101110111111010110100110011001010011011110110100011010100111101001100100010101001111001100;
    #100 Din = 128'b11110010011101111000010001111100011001011101000011000100001000111100100101111110011011100110110000001001001000010101011101111000;
    #100 Din = 128'b01000000011000101011110111100111111111010110100011100101111100101101100010110010011001111010101010011111110001001000111101010011;
    #100 Din = 128'b10000100101001110110011100101111100101110001011101110011110001100000110001010010111001011100000100101111001101011100110101011001;
    #100 Din = 128'b11100110010000100000110000010010111001010001101110001001010110110101101000011110000010010100101101011010100001100101001110011110;
    #100 Din = 128'b01110010000101001101000001011011011010010000000011010001100001011111011000011101100101100001011100110000010101111000001101110011;
    #100 Din = 128'b10110100101100101101110100111111100111000111000000110000010101011010001100001011100000101111010100001011100111101010111111100011;
    #100 Din = 128'b01110101001010110000110010110100001111100000001001110010000010010011011111110110111011000001101001000111011110110101001000000011;
    #100 Din = 128'b11110100001011001110010101001111011110111001111110110110111100101001100111101100011011010110010000001101001000111100101110111011;
    #100 Din = 128'b01101100111000001000010011000111100110101101110011011001111010110010001100110101011100011111100111110000101101100101011010001100;
    #100 Din = 128'b11100100001111000011000001101100110101000010011011110110001111000111100111101100011111111010001001010001000011011000011010000011;
    #100 Din = 128'b10111000001000100001001101001001100101001111000001101011001011101001101100011111011011110001010001001110110100100011111000110110;
    #100 Din = 128'b00100000110000000010111000000101011101101011100000001011000000011110010001110001011101101100011010111010110110000000100001010110;
    #100 Din = 128'b00010000000011011011000110101011110000011001100101101101110000101011010110010010011010001111110111110010100010001000010101010010;
    #100 Din = 128'b10110110011111111111000010011100111101000001001101111010100100101001100011100000011101100000001111110100000101001100011011011001;
    #100 Din = 128'b01000110100100111001001111001101001101110011100101111010110101110101100110110101101001111110001110101000100010110101101000111101;
    #100 Din = 128'b00001010000101011101000011011111001000110010101110010010011010011110010111100001010100100010011111001110010010010101000011101011;
    #100 Din = 128'b10011110011001000101000100010001111010001001111010100101110001101011010010011110111001000101010110100110111110111100100001011110;
    #100 Din = 128'b01101011011001000100101111101100001110110101101011100010011000100000111000011111001110100111110101001100111011101101011101111100;
    #100 Din = 128'b10111101010101111011111111011100111000111110111011101110001101010100001110000001110001110110101000011110110011111100001001011110;
    #100 Din = 128'b11101001000111111100010000011111000011001111111101110110001011000101100010111001011010111111111010100111101101010000111011010110;
    #100 Din = 128'b01000111001100000000000100000000110000011111110111110100010010111111000001100010110000101010001001000000011001101001101011111000;
    #100 Din = 128'b00000100011101100000001101110101000011110101100111101010111110000011000110000111100001011101111101000000101110111011100001011001;
    #100 Din = 128'b10101000111001111000101011110011011110100101110111001100100011101010110101110010101010000110110101011010111011001111111010000111;
    #100 Din = 128'b00100001110100110010111010010010100100000010110000010000001110010110100011100010000011111001000101101011011001101100010101110000;
    #100 Din = 128'b00011111001100110010111010010001100100110101110111011000001100111011111100000100000000101110111011011101010111001011011001011110;
    #100 Din = 128'b11010101111100110100001001000001000110000001110101001010110101100100111011110111000100001101010100000001001101011101011001001101;
    #100 Din = 128'b00101101010110000110111110101100101100101100011001101101100100011001000001111001010101111100010111110010000110100111100111100101;
    #100 Din = 128'b10110100111011110110110100100100000110011101011001101010100111101111011100100010011001110001100010101111000001010010100101110010;
    #100 Din = 128'b11101100101011101100111011001011000100010010110111011111111000011011010111110101010111100011000011101000011111111011110100010001;
    #100 Din = 128'b01010110001111000010101111101011101011000101010001010001001100000110100011111111000010010101010011111001100110010011111011101011;
    #100 Din = 128'b01101010110111010000100011010110000011010100110001010100111110110010100100110111101111110101010010001000110110001100110001101000;
    #100 Din = 128'b11001111011011000100110000100101000110101100101001011101011010010000010110111110000000101000101011101001011100000101100100110011;
    #100 Din = 128'b00010101111110101100101011001101011100010000000000010111010001101001111011101000001011110000011100000001111000010100010011101111;
    #100 Din = 128'b00010000111011011001001011010110001101111000011010011100101000100011111001101111100110010101111101010001001000101001100111000011;
    #100 Din = 128'b00110101001101110111001011111001111100111001101110110110101101000100111100010101010011100111001110100110100101111101011100011101;
    #100 Din = 128'b00111100111110000101100010101010000001001001000011110101100001011010010010000001000100101001100001001011111011000111011000000100;
    #100 Din = 128'b00010011000010010111011110110100100100010001011111010100010111100101000001111110100011111001011111111010000001111011111100101011;
    #100 Din = 128'b00011100000100011101011100011001100001000101000010111011100010000110000011101010011011001010001110011100110100110001100110001010;
  end

endmodule
