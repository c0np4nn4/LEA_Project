module LEA_EncDecEXAMPLE_tb;

wire [127:0] Decrypted;
wire [127:0] Encrypted;
reg [191:0] KeyIn;
reg [127:0] TextIn;

LEA_EncDecEXAMPLE
 U0 (
  .Decrypted(Decrypted),
  .Encrypted(Encrypted),
  .KeyIn(KeyIn),
  .TextIn(TextIn));

  initial
  begin
    KeyIn = 192'b010010000000100101011100000100010110110001010111110111110100101111100111100111110010100110000100011100001101010011000001010010011100011110111100000110111101101001001000111010011001000011010010;
    #100 KeyIn = 192'b011011100001111101001101000000000101110011101110011001111010010100010111001000100010010000101111001100000001110100001011001000011001100111111111111000010110110100110111010101111100100011011001;
    #100 KeyIn = 192'b011100011001111100110011000110110001110010000011000110010001100001011101100011010010111010100011000001110010000110101110111011001111010000111110000100011100011100111111001010100010111010100001;
    #100 KeyIn = 192'b000010101001010101101010001011000000000110111001101101001101110100011000010110111010111111111001011011100010111100011011100010000000000010010000100110100011101000110010011101110111001110001001;
    #100 KeyIn = 192'b110001000010101001101011001011111011000000100100001000100111011100010000110010111010100110011000011011011011110001110010001010101111000011101011001011001001011001100101110001000101111101100000;
    #100 KeyIn = 192'b111011001011010110010110011100111001100110010011100101001010000010111010101001100011110001011111100000100010111111100001001110011110110010001110011100000010100001110010110110101000110011111010;
    #100 KeyIn = 192'b111010101100011101001001001000001001100000111100100110111000000111100100001001100101010000110010100101001000000101111101110111001010111001001101100111010111011000110001010010010100000100111011;
    #100 KeyIn = 192'b110000111001000010110101100011101000011100011110100101001111010011011111010010111100110111000110111100110001110001010101011100010101110100110010010000011001101100101101001110111101011100010110;
    #100 KeyIn = 192'b011100101001000011000111111010011101010011100100111100001110100010011110010100001000011010111101010100111100001000100110101010110101110100111100010011100101110001010001011101101001100001111011;
    #100 KeyIn = 192'b011001010001000001011011100100001000000000101010001101011110011000010110111110011011001010111011100110101111011010011110001111011111000001010010111101111001110101100011010111111001101111011101;
    #100 KeyIn = 192'b000100111010110110111111110011001101000100110000000010101111011100100100000001001000010000111001100011001001001100010000100101110100000100010101110110101100001011111001110000011101110011011101;
    #100 KeyIn = 192'b101100010111100101000111001110001111110011010000011101010000001001000001010101010011111111111001100001010001000100100011010001101001011110010101001111100001100011101010101000110110011000100111;
    #100 KeyIn = 192'b001111010000011100011011000011011110010011011100011111101011110011000100010101111111001110000001101101110001101101000100001111111110110000010001101100101011100111000110010110110100010001110000;
    #100 KeyIn = 192'b001000111000011010101010101001010101001111110111011100011011101000000100111011010000110000010000110110100001101111110000001100100010001010100011110001000101100100010111111000010011111010011000;
    #100 KeyIn = 192'b011001010100111011001010010100010101100110101110101111010100011001111011011111111011010110111101111010100010010111101001011110111011100011111101110100010101000100000000100111111001100011000010;
    #100 KeyIn = 192'b110110001101011010110011010110011111111000100101110010000000011111000011011010111101010010110000011101111110111111011000110111100000001011100111000101111111000111001111010110000000100011010100;
    #100 KeyIn = 192'b010000100011110110001101001100111111010110110010010010011111010110000010000100011100110001100111110000010100101001100000011000011010001111110011011110101111100001101010101001110011100100011010;
    #100 KeyIn = 192'b001001101101111111000011010111100110101011011011001010111101101011111101101101111111110100100000101100001101001111100111000100011111001000101100011111011101111110101101011100110000100010100111;
    #100 KeyIn = 192'b110110101011100001000010011110000000101100111011111001100011011011011011000010110001110010011010110101100111101111000000011101110011101001000000111001110101001111110010100101000111010010011110;
    #100 KeyIn = 192'b000001010100101001110000011101110101101100000000010001000011111001110010001111111001101000101100000011100000011011110100011001111001000100010011010101000110101111100010110000001110101100010110;
    #100 KeyIn = 192'b010110100110111001001101101000101010000100100011110111100010101010000011100100101000010111010001100010101101001001101100101001110001110100111101011001011101011111010100010001000001011001010011;
    #100 KeyIn = 192'b100100010010011101110101111111101010100100000001101000100011001011110001110000111111000110100000111010111010101000100000001110110110100101010000011011011111111111001111111111100001010101011010;
    #100 KeyIn = 192'b010010100110001001011100001100010011001101110010101011001000000101110011011001111110000001010101010110000101001101101101110010100001000111011110111001100111000110000011000100011111000100110111;
    #100 KeyIn = 192'b110100000011011111101010001001011111010101100010001101001010101111111001111100110001010000010000111100100000011010001000000000100000010010010101000001011111010010000000010010100001010000101110;
    #100 KeyIn = 192'b101101111110011110100010001000001111111010110101100100111110100010110000000100011001111011110110100111100010011110010100010110001110000100101101000000101010110110000100001101010010011101110000;
    #100 KeyIn = 192'b011110100001101111001010100001110010000101111100001111101111011011011001110111100011111110101100001110001110001101011011010111100000011001110100000101001000010000001010001011011000101110111101;
    #100 KeyIn = 192'b010100000000111000011111011000010111101011011011001101100100000000010010100100110101100110011011011000100111101010110110100101100110000111111000100110110110011110100001110100101010101101101111;
    #100 KeyIn = 192'b011100010100011011011000011111111000001100010000101011101111111101111111100011001100000010101111000100001101110101000100111011101001100111010101111101011010011011101101100110100000000010000110;
    #100 KeyIn = 192'b110000110110110011000111000100101111110101010001111010111111110001101010001000100000000000111010111010110010101101000010101110100001010001001010010100100000111111011001010010001010100101001110;
    #100 KeyIn = 192'b111010000110010110110101111001101000111011100110100011111110011111111000100011101111101111111101001000000111101000001110000000000010001010111101100001101110101101000110111100001110001001011011;
    #100 KeyIn = 192'b101001111111010100111000110000100000001111011100101101010111100111110011010001000001110001100101100000001000000100010101011111000010101111011011111011010000001011101101100101001101001011010010;
    #100 KeyIn = 192'b111101110001100001010010110101110111011101000010000000111101111101100100100010100000011100011000111011000000011011111011111000000011000110110101100100010011111110011011000110000001101110110101;
    #100 KeyIn = 192'b101100001101000011011011100110000110010111000000000000110101011100101111011110101011001110000010101000000101111010111101001000010110001110101101010011010011100001100000010010101010110101111111;
    #100 KeyIn = 192'b111011000011110000000101100011011110011011100010110010011011101001011011111101110101110111110011000001111111100110000000010011010011111000100011111001001011101000011111111000100110010100001010;
    #100 KeyIn = 192'b010010111110000101000011011110110010010010100010110001110100000110010011011010011011000011010011010111110100001000010111001110111001110110110000100110111101100111100010101100001111111100000011;
    #100 KeyIn = 192'b101000010010101000010010111001001111000000100101100110001111010100010001011100000000001100010000011111010010001010100001011110011000110100111000111001001000100100111001110011101110100010110111;
    #100 KeyIn = 192'b110011101001100000010010011100101100111010011101111001010000100010010100011000001100100011001010000101110110100010110101011100110001100000001110011001011001000001000100111101001110101111010101;
    #100 KeyIn = 192'b000101010011000111001001010111111000100101111011010011101000101001011010011001110010000011111000001110000001100101000100101010001111011111001101010000000011001101100000001101001101101001100110;
    #100 KeyIn = 192'b010011110101001011011100101100110000100110100000100100100001100010111000001011000110101110101001101010010011111001101111001010111101010101001000011100110000101110111110100100011110100001111101;
    #100 KeyIn = 192'b001111101100001111110101010011010111100110001011100101101101111010110110010110110100110001110011110001101001001000010010001101100100111110111000111100001000000010101001011111001001001111100011;
    #100 KeyIn = 192'b110011000101101011001010010000100000110101100100011111101100000101010000111010010101000001010100001010111110011011110010011111010110011011011000011100111110000111111101001000001110000101000110;
    #100 KeyIn = 192'b111001110011101101000011001010001000101110110111100000100010000010100110001001011011000100000011111100011000101001000100010110100110100001011110111100011110010001010010110010111110001001100001;
    #100 KeyIn = 192'b011101001001001111100111000111111101101011110111110110000110111110001001001000100011000110001101011100001010011011101110011010011101101011101010110001011011000011111010000100111111110010010010;
    #100 KeyIn = 192'b100101111011110111010100010010000110101000100100110011110100001000010010000011110111010000000011001110010100111101101101101100111110101010011111010011110010011100100001100100100100111001110110;
    #100 KeyIn = 192'b111111111110101100011110001101000100010010110100000010101110100011000100101001001111110101101000100011001011011110010110100000011011110111011101110100110101100111100010001111101001010100110101;
    #100 KeyIn = 192'b110111101010100101111101000101000101010101101011001010101111100111000000011000000010010101001110000111010111000101111100010111100110100001011111000111000011100010001001011000001100011011000000;
    #100 KeyIn = 192'b101001001101011001001101100010010110100011000001011001010001111011000111110010101100101010100111001101101110100100101001001011110010001000111100011010011011011001111001010011011111000011111011;
    #100 KeyIn = 192'b101011110101111011111011101011000000100111010100011010010100001011010010101001110101010010011110001001010100000110010011010000001111100001000101110100110110111011111110111011011110011110111011;
    #100 KeyIn = 192'b010000001001110100011111100101011100111110101101000110000011000111101000011101101101000110110100000000010011111110010100110100101110011011010000001100001001011111100100111101101101010010101110;
    #100 KeyIn = 192'b000000111010101111000001001000110100001111010111010110100100010100100000001111110000000111011110001010111000111110110000000010111110010101111100100111001001100101010101010011101111110111000000;
    #100 KeyIn = 192'b100110101001100101011010011000110100111000001101111110000111010000110101100011001010111100111111100101111110010111100111100010001100011101010000011100111100100100111100010011001010010101101110;
    #100 KeyIn = 192'b010111111011001011100111011011100011010101101011111000111011011110101010011011001010100100100101001110100011110011110011010000111010110001110010010101010100010100101011010011000110001000001101;
    #100 KeyIn = 192'b100100100001000000000010100101001110100100000011111010010000001110110100011110011011001000100010110011001010001110110001000101100001011011111100010101111011101110011001001010010111001010110000;
    #100 KeyIn = 192'b100011110010001011110111100001101000101100100101000010111000100111011101001110101110011101110010100111001111011111001000011111001111011000010111001101101000111001101011100100011111001110101010;
    #100 KeyIn = 192'b000100101101111111010011011110010001000111110011011110000010101011011111011011001001111001000110101001000010000101010011000011111111001110011001001110101110100000010100100000010110000000100001;
    #100 KeyIn = 192'b110010111100011011101110110111001001100100010111101101011000001111100111010111011101010000000101100101101000110011111101000010001000001010011001110100101110101010010010010010111001101001100010;
    #100 KeyIn = 192'b000000101010100110001010110010111100101110100000101010011101110111000010001010101100110101100001101101100111111011011010010011111011110000110010000100000001111110101101000100100100010010110100;
    #100 KeyIn = 192'b010010110101000110101101001010110010001110100111101011001101011110100111100111000110010001111111000111100010100011110111001111101101110000111010001100101100100010101101000011000110110010101011;
    #100 KeyIn = 192'b111110100000001010101100111001101011100000000010000100101001111000000101001111001111010111110100010001110001001000001110100100110001111110011110101100010000100100111111000000001111100011000100;
    #100 KeyIn = 192'b101001000100001110101010000101000001111111010111111101011011001011111010101101001011101001111001000010110011000101000111011011111101111000101010111011010110001101111110011001111010100111101100;
    #100 KeyIn = 192'b110111000001111110000000110011000001100001110000111011111110000011010001000100110101001111101101000000000111101011110111100001110000100001111100000000001010010110110000010101101101100101101001;
    #100 KeyIn = 192'b100011001000100101101100010100110101101110010001110111010000100101010001101110000100000001011001100010011101011010000010101010100000000101000110100000110011100000010010001101011011011010111010;
    #100 KeyIn = 192'b110010001001010011110110110100011010011110111100011100010001111101100011101010001101111011000011110010101111101011101001001000101110010001110010001010011110011101010001000010001011101111111000;
    #100 KeyIn = 192'b011000011111111110100101000000100001000011000111000100001111000011001111010100001010010001110100110100100011000111001001010111100100111101110010100000101101100000111001110011101111111010000110;
    #100 KeyIn = 192'b011101011010110001001000111100010100100111110000001000111100011100110111010111100010010101001111100110100111111110010101100110101010100010010011110011101000100110100010000110000000100110010101;
    #100 KeyIn = 192'b101010010100001011110010011101110000100100101101001110001010000011010100001110111011100111001100110110001011010111100101001000100101100110011000111111000010110001100100100001110001101011001001;
    #100 KeyIn = 192'b111010011000110111100000111001000000001010000100001001100100110100111011100011110100101100011101010111001011111010101101101011110011011111001101101100001101100001000000111010100011100100100001;
    #100 KeyIn = 192'b110111111101001001010000100111100110010111000110110100111111001111000000010010000101100001011111111000011111111110110100110101100111111101100101011000100000010001100111111101001010101001001101;
    #100 KeyIn = 192'b000110011011110000000011100110001110001110100110101001110111111110011010101001100001001000000100111110100111100010100000111010010000101110101101010010011010110101010000001100100111101101001100;
    #100 KeyIn = 192'b101000100001010010101000100111100111100000101100001011010100000111101011001000100000010000100111011000000110010010000011011101011101100001001011001011011101011011011110100011011011101101101110;
    #100 KeyIn = 192'b011110101011111110000101111100111100100000110001011101111111111000001110011011011101011010011011010011110111111010000101100000010111100100111101011001011111110101011111001011101000101010111000;
    #100 KeyIn = 192'b011001010111000110101101011110011100010001110010000101001010101001000111001000001001011000011100011101000101010100100110111011001001101101011111011001101000111100101000100100010011010100000000;
    #100 KeyIn = 192'b101100000110111001101011010101110011010011010000001101010010011011100010100100011111110000100001011000000111110110010011110100011111111000101100100100110001001000011100100010000101001101101101;
    #100 KeyIn = 192'b100000100000011010100010000111110100111110011000111100110100110000011010110111111110000101010010010111110100110100001001110000101001001110010001011001010111110011100110000010100000011111100001;
    #100 KeyIn = 192'b010100011111111101110001110100110111100100111110000111111001011111000011110011101100111000100110011011011010000011010100010011011001100111010011011101100001100111110000110100100001101101011110;
    #100 KeyIn = 192'b011011101001100101110100000111100000001000001011100111011010111100000100000010100011111011010110110000010011100010011010000001001001010010101011101100010011111110110101110101001101101110110101;
    #100 KeyIn = 192'b001001010100110011011011001000001001000010010000001110111100000001001011101101000101100111011011111111010010101110111000000101011111110001000011101110011111101101010110101010010101000000000000;
    #100 KeyIn = 192'b000010100010110111100101001000000001000011001000000010001111111010011010011110010000010100111110100111001101001100110010000100001011100110100000010111111110011010101011010110001101101100101101;
    #100 KeyIn = 192'b101101100110110011011111101011101010011110100000100001001010111000111011111000101101010010011001010100110100111000010001000111110001010110001000100010010011001001100110111110101110110000000101;
    #100 KeyIn = 192'b010010011001111001101011000010110111011000110101001110010111110011100000110001110000011100110111001011100111010110010111101000000010111010000110100100100100011100011000110101110011000001101011;
    #100 KeyIn = 192'b010010101111000101111000111100001100111000011101111110011100111111011101101110100001001001010001101010000000011101111011101000010011101111111011101110001001010000000000010010101100011000010111;
    #100 KeyIn = 192'b000101101110000011100101001100010011000100111111011000110101000101000101110010011111011010111101100100000100010001000100001000101010101111001100111011100001011111110000101110101010111110100000;
    #100 KeyIn = 192'b111010000110110110100001100110100100100100110010000001011100000000101100110001101001010100110001000011000101110010011010001111000000011001010101010010100110011011000110100010100000000010010001;
    #100 KeyIn = 192'b001000111100100110101010111110101001111001100111101101101101111001110101010010011000101100101101110010011010111010110000011110100010000000101100101111111011101011101101100110111110111101101111;
    #100 KeyIn = 192'b000010101110100111111000011000001011100100111010010010010011001010111110000110110110110000010011010001110101011010100011010101100110001011000111000100001001110110101000001100101111001001111101;
    #100 KeyIn = 192'b101010000100001111011011101111100000010111011111110101101110000101100111111000000011101110100101110001001100100111010111110011101100011001010000000110111111101000100111100000010111011101111100;
    #100 KeyIn = 192'b010111111101000110001010100001111101110101000001111111011001101000000111010100111111110011101100011100111101010000010011000010110110100101010000010001000101011010011110001010110010011111010010;
    #100 KeyIn = 192'b101100000011011111001111010101011111111000110110001001111101101010001111110001111010111100101001001010100100010110001111001010100001010000011111100011111001011011011101100110001010101101011001;
    #100 KeyIn = 192'b111101001111000100100001010100001011010000010010101101001110010011111111101110101100011011000101010101010011110100010000111100101111011111001110101010011100111000010001110100111000010010101011;
    #100 KeyIn = 192'b001111100110100010000000110011011100010110011100010100011000101001011110000110001000110001111110010101110110010010011000101101111101011110010101000110111101101011001100001111011010001101010010;
    #100 KeyIn = 192'b101011010010010100110010111010111011110011011000111000000110000101101010111110100010111100101111110010011001010000110010000100100001110011010011110111001100001110111000110011111011001000001110;
    #100 KeyIn = 192'b011100000100111111100001110000101010010011000010001111011011011110000101100101001111100110111000101110100101010011010010101001010010000000000110110000001000111001001100100000011111001100111111;
    #100 KeyIn = 192'b010011100110000001101111000100011011100011000111101011110011101111110110001010101000100001101110110010010000001101011011101001001111001111011111111000110101000001100110101101000011110010100010;
    #100 KeyIn = 192'b111100001100110011001011111001101001000011001100011100000101001100010001001111100000101000010110011000001100101011110100011010101110000000111100110001011001000000100101111100100000110011000000;
    #100 KeyIn = 192'b001110110011001111111110000110000000111011010110110001001010111101001000001111011100010100000111010100001111010110100010100101110001010110000010111010001011111110010111111011111101111100111101;
    #100 KeyIn = 192'b101001011111010011111000001011011110110111001110111001001000000111110100111010011010011001101001011011011000011000110111010111110110100100110010100001100010010101000001001010001110100011111001;
    #100 KeyIn = 192'b100000000100100100010100000001100011010001110000111111011010000010000010100110100000010101101000100001011111000011101111011000001010100011000110000111101001011100001010000111110110111101111000;
    #100 KeyIn = 192'b110111011100111010011011010001010101000110100101111111000010110001110111111100011100111010001111010011100111011101101110111100111101101000101100011010010000111101000011110100101001011100001101;
    #100 KeyIn = 192'b011000011101111100010011010111111001111110101001000110011111011101000111000001100010010110000010011101111111000100011000100100100011100001000100110000100011011110111100001111011101010001110000;
    #100 KeyIn = 192'b100100100110010011110000110111100101010100011111101001110010101101100110001101101111100001001101001101110110110010000010111101011101000101101011000111100000001010111011100000011010001100010010;
  end

  initial
  begin
    TextIn = 128'b01001001101100000001001000110111100111101111000001001111101111100011101000001100000111111010010010001001111110010011110101000000;
    #100 TextIn = 128'b10110011010010111111100001100011100001100000001011010010011011110010101010110101100100101011000001100100100000100111011110010011;
    #100 TextIn = 128'b10101001101011001101000000000110111111010111101111101110100101111111101100101010010011010101000100100011110100001010110100100010;
    #100 TextIn = 128'b11101000000110011100110010101010011010111000100101000110110110000111011101010110111101111101011001010110110000000001000110111110;
    #100 TextIn = 128'b01100000101001010010101011010011101001010110000100110101000001101111100000101001010011000100100100011011011001110110011011011001;
    #100 TextIn = 128'b01100000010001100101000011100010001101111000011100101000110000011000011111011101111011000100101111000111101101001110101000000110;
    #100 TextIn = 128'b10001101100010111010100110000100001000111011010001110101101111100000101011000000110100100011101000011000100001001101101111110101;
    #100 TextIn = 128'b11111010010011010011001000001101101000110000101000010000100001110000010000000000111110101111100110111111001011011000000011010101;
    #100 TextIn = 128'b01001100000010000011100110110010100110110001010010011010011011100101111100011010001001100110011110110000111111100101011011011110;
    #100 TextIn = 128'b10100011011000010110001111111110010101001100000100010111101001101000111110001111010110000000111001010010111010101010001000110001;
    #100 TextIn = 128'b10000111001101100000001011011001110010101001011000110001011001111000101010011011110110001100000100101011111101100001111110100001;
    #100 TextIn = 128'b10111101111101001110010000111011010110001000101110111100001010011000110010100010010111001011000001011011010101000001000001101100;
    #100 TextIn = 128'b00000111001101010000011011010010010111010001101001000101010111000100111000000011110011110110000010101100100000100001101110010101;
    #100 TextIn = 128'b10001000001000101100000111000000000011010101100110001001101011001101001010101111011100110101101100100011011110011000110000001111;
    #100 TextIn = 128'b00111110111100000101110001111010000100001000110010000101101101100001110110011011011101110111011100000000011111110111100110101111;
    #100 TextIn = 128'b11011011011001100101110110101100010101111111101001000001011011010010110001111010111000100101000101011001111011111101110110000001;
    #100 TextIn = 128'b01101000101011001100001000101100010000011011101000101000110101100100100011010011111011100000011011010101011010010101101001101100;
    #100 TextIn = 128'b10110100000000001001111101000000111110010001110100011000110111010000101101100101001010001110101111011110110000110011110111111101;
    #100 TextIn = 128'b10100010010100000110011101001101100001010011011110000110011100110001000001111000111001000111100101000100111111000000110000111111;
    #100 TextIn = 128'b10101100011010001101100101000000111100110001111001000011000100011000000000101000110011101100010110101101001100010101001000111000;
    #100 TextIn = 128'b10110010111111101011000010011001011011000101011010101100101001111100101011011011100101101000001101101101000000111000011000011010;
    #100 TextIn = 128'b10001010011000101100000001101000101110010011110001011010001110001001001001000101001100101101000101110001100000011011111101101011;
    #100 TextIn = 128'b11010111111000011011101110000010010011010101101110010001110001100100100001111111101011100011101111101101110110000000010110101100;
    #100 TextIn = 128'b01101010000011111001000000011111100101000000001010010000101101110110111001000101000101100010101101000011110100100110101111000010;
    #100 TextIn = 128'b10110111111100000011001110111110100001010101110100011110011010010011111001110001101001110111011000100101010110100111010101110110;
    #100 TextIn = 128'b10001101010110100010100101001101011100111110100100001110010000011000000101001011000111110011100000001011110000110001011100000010;
    #100 TextIn = 128'b01111000000101111011010110001101101101001100100110011011101100110010110100110000001010101101100101110000111010111000001110001101;
    #100 TextIn = 128'b00000010011001111111101101000110000001101100001000101001111110000111011100111011100110011100000000001000101100010000111000111000;
    #100 TextIn = 128'b10101101000010101001001100100100010001011100011011011000001101100010110010000010111000000100100100110010110001100011001010110100;
    #100 TextIn = 128'b00011010101001000111101110000101111001110000100100000000110100110100101100011110111111000111110010100100100011011110111111101111;
    #100 TextIn = 128'b10110000101110001100100001100100001011000110010111001011011000001001000010000100110111111111110111101000100100001101101101111101;
    #100 TextIn = 128'b10010010110011101010000011001101110110110111001111010111000111011010110011100101001001111010110101111111111011010011101101010110;
    #100 TextIn = 128'b11001011010110110101111111011100010001111011101010110010011011111010101110010111110110100111000010011001010010011101010011011101;
    #100 TextIn = 128'b11010000101000110001101010000110011011000010100110111000010001011011011010111010100101011010011000001001010100001100110101001111;
    #100 TextIn = 128'b01010110110100011110010111000111101000010001101001001000001111000001110011001111000111100100000000110111010110011001111110000001;
    #100 TextIn = 128'b01100011001100001000001100110100110111000101110111110001110011010001110111101100010010001001100011001100001010001010000010011111;
    #100 TextIn = 128'b00010001000001110010100010111100010100001110100010101001110100111010110100011110110100010100000001010011010101111011011101001000;
    #100 TextIn = 128'b11011000011001100010011101000001100100101100111101010000010110011000010010101001010010010001111011100001110010110011010000001011;
    #100 TextIn = 128'b00001010100010000011100101011010111111001010101101010011001110100110001001001111111111101001000011111010101110111110011111111111;
    #100 TextIn = 128'b01010011111001000110011001001001110100111000100111010100001110100110101110110111001101010111101000101100101000000101100010111100;
    #100 TextIn = 128'b00000101111111101011101010000010111011010101011001111110100001001011110000111110000010010100100101110011111111101100001011000110;
    #100 TextIn = 128'b00111011010100100011100101011011011001111011011000001100011000110010110111111001110010110001110001010001110000001110111111000010;
    #100 TextIn = 128'b00110000101101001111011110010111010100111000101011110001010100100110000010110001101100100111111111010110001001010100101001100011;
    #100 TextIn = 128'b01011110010111010111010001000001011111111100101011111001100010100100110110010111011011110100111101011101010110000100011111001111;
    #100 TextIn = 128'b00011100110000011000101001011110001111111011011111101111010101001000100100111001000111001010010100010110000101100000010000010100;
    #100 TextIn = 128'b01011011100101001101110010101001000111101010100100010100000000111111100110000100011011111101011010010010100010011010001011111000;
    #100 TextIn = 128'b10010001100110000110001101101110010110111100000111111010011111000111010111011001101000010001010011110100100011000001000011111010;
    #100 TextIn = 128'b00010110010100010101001110001001110001110111000011101101101011001000111000100001101111001000010101000111001111110100010101011011;
    #100 TextIn = 128'b00100011110100011100100111101111110010011101010000010101001010100010111001100110100111011111001011011101100010011110110110100011;
    #100 TextIn = 128'b00110111111011010101100110100100101100100000101001101010000011000111111111111110100110111010111111110011110110111101100011011010;
    #100 TextIn = 128'b00110111101011011010011001000110111000000001000011001010101100000011111010000001000111000100111110001010010000111110111011001011;
    #100 TextIn = 128'b01101111110111100001011101100101100000010001111111101010110011111011001010011101011001101010010010011010110100011011010000100000;
    #100 TextIn = 128'b11011001010001000001011011011010111100111101001101100101101100010100110100011000100001001000111101000011110001111111010000101010;
    #100 TextIn = 128'b11101001100111001000001101010010101111111110000110010110111001110100011101110011111100001001010111110100011011110111110100011101;
    #100 TextIn = 128'b10111011100111101001101001110011111110010000010110100110111010111010110110111000101000011011001011010111100110111000101010011001;
    #100 TextIn = 128'b01011011001001101101000000110101001111000110100111111011010000011101011011001000100101100010010100001100100000101010000000001001;
    #100 TextIn = 128'b10000100111100110010001011100101110011101101001111101100111000101000010110011001011111100010100000111111101001101011101001001100;
    #100 TextIn = 128'b10101100110111010111010101000011100010010011101000011010100001000101001111100011001001111001111001010000111011111101011011000010;
    #100 TextIn = 128'b11100000011010101111101110101010010101100101000111000000010000011011110110010000011001111000010101000010101011011001110001101111;
    #100 TextIn = 128'b10101010011011001010111100000111111010001100000011110000001100001100010111011010111011110001001000101010010100100000110111000100;
    #100 TextIn = 128'b10000100000110101010101110111110011000100011111100110000001010011001010100011110101100011001111100101101000110100011110111110010;
    #100 TextIn = 128'b00011111101111001010011010111110110111000110010100000001000101111011011101100000100100001111010011010001110110011100001100111110;
    #100 TextIn = 128'b00111010001011111011010001010000011110011011111001011010101000100111111101101001000011001100000101110111111000110010000100001001;
    #100 TextIn = 128'b00100110100101001111011100110011001010101001101001101000110010111011101000010011110000011001111010101110000011011010010110101111;
    #100 TextIn = 128'b00110011100011111111000001011100101001110001100000110001000100000111000010111111010110011110001111011010101101011111111011000001;
    #100 TextIn = 128'b11101001011001110000100000100011010111010010111011011111111111101011011100101101001000010100100101011101110010000110110011011001;
    #100 TextIn = 128'b10011001100110100011010111101111000001101100000001010011010100000110011011011000111111011101011110001010100101100010100110010100;
    #100 TextIn = 128'b10010001001011100000001100111101010100110100101001111101011100110100001011110000101101101000111100111010010011011111011011110111;
    #100 TextIn = 128'b00010001010110110000111000001000011011001001100101101000110001101001010101000111000101100110011100110011000111111100010010001100;
    #100 TextIn = 128'b10110011101100010011011101000000010100010000011000010011110010100001101000000110100011010101010110001110101001110100101010111110;
    #100 TextIn = 128'b01101100011000111100111010011100000001010010101010011101110011000001101101000000011010010111010101011100101000000111101010011101;
    #100 TextIn = 128'b00000101111100111011101111010101000101110101110111001010100110010001001110001110001000110000111111000000001001000000010000110010;
    #100 TextIn = 128'b01011110001000011101010010101000011110100100010010110110101010010100100100011011111100011101000101101000101110100010101111011100;
    #100 TextIn = 128'b01101001010001000111011110011000101101111111010100001100111011001011011000001101111100011001100001000110011111000011111110100010;
    #100 TextIn = 128'b01010100000011001110101101000111011111101010000010101011100000111001101001110101010111110111010011001011110001101100011111000010;
    #100 TextIn = 128'b10011100010110000011001010001010011110010111010000100100001000011001001011010001000011111001001101111010011010110111000010100110;
    #100 TextIn = 128'b10011010100000111111010100110010011110101110111010011101010011101011101100111001000100000001011001100001101000100000011011100111;
    #100 TextIn = 128'b00110100000110010001000101111011000010001100110101100110101000101010100111110000000000010011000100011000110110001111100011011010;
    #100 TextIn = 128'b11111101101001000010000010100000110111011101101111101110101110110110011100111101001011001110101111111101111100111101100010011000;
    #100 TextIn = 128'b10101111110100110001000000101111111001010000110100001000000110011111000001011101000010101101000101001110001110100101110010010101;
    #100 TextIn = 128'b10110011110110010011101100001001110000111010001010010000011101001001000000011000101001011001101111010101011110010011011011111101;
    #100 TextIn = 128'b00101010111101111001110100011110100000011110110010001100101100000110000011110101001101111100111010011100101000110110100100111001;
    #100 TextIn = 128'b00000000100111000010000011110110101100010111010011001100010011010010100110101000011001011001001011001110011011000101111101111110;
    #100 TextIn = 128'b11111010000101001101001110001100010011001011010101100100010101100010011010010111101110001101000110001011010011001010001000011011;
    #100 TextIn = 128'b01011110110101001111111111011111000110101111111001110000111101110001010101001101011010101001010101000010001000111000000110011101;
    #100 TextIn = 128'b10100100100011001101110111111010010101100110000110100111010001011011001111100010101001100011110110100011100000110001011110001011;
    #100 TextIn = 128'b11100101011010010100101111110110111111101010100011111101011110001001000001110010101000100000010000011011010101000010001101000010;
    #100 TextIn = 128'b00010110001011110100011001011010100001111100000001110101010011111110011110111111110110001110110011111001101011101100000111110000;
    #100 TextIn = 128'b00010001001000010100110010111000001010000011010100000001101100100000101001110001010100101001100110001010110001100110011001000001;
    #100 TextIn = 128'b01111010010010110010101001010010101001111111010010101010001010101000001110101111000011110111011001101110001001110111001110000101;
    #100 TextIn = 128'b10000100010000001110001100111111100010111011011101100111111010100011101000010110100111100101000010011111100000111111110101001011;
    #100 TextIn = 128'b00111101111101011111111100010101101000101000000000011011100111000001101100111110111100101010010101000101111110100110110110001000;
    #100 TextIn = 128'b11001001010011001100000110111001110111111110001000111111011100010011111011000000101011010110110011000010001010101010111101111010;
    #100 TextIn = 128'b10111001011101110111011011010001110000011011100001100000001001011010000100101001111010101111001110111100000000001100100000011110;
    #100 TextIn = 128'b11101110001001110010001000111111001100100001001110110110001101110100110101100001100101111011110111110110010100101110110101101010;
    #100 TextIn = 128'b11000001000010111010101010011110101101101101010011000001010111011100001110111011000110010101001101001110001001000000010101101010;
    #100 TextIn = 128'b10100100011100101001000010010001011000011101101011101101011001110111010001000000001100001011100110110100000011010111000110010100;
    #100 TextIn = 128'b00011101001110111110110110011010110010111111010110101001111101000101100000011010100110000110101110011100001001001100101111101001;
    #100 TextIn = 128'b01000000000000111110001010001111000001100000000010011011100010101111001111100101000111000010101110000011101010010101100000111111;
    #100 TextIn = 128'b00010110011110001101111010000010110001011010001010000111010100110001010000000111101101001001011101110001110011010111001111110110;
  end

endmodule
