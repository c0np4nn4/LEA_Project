module LEA_BlockSubtractor_tb;

reg [31:0] A;
reg [31:0] B;
wire [31:0] Result;

LEA_BlockSubtractor
 U0 (
  .A(A),
  .B(B),
  .Result(Result));

  initial
  begin
    A = 32'b01001000000010010101110000010001;
    #100 A = 32'b01101100010101111101111101001011;
    #100 A = 32'b11100111100111110010100110000100;
    #100 A = 32'b01110000110101001100000101001001;
    #100 A = 32'b11000111101111000001101111011010;
    #100 A = 32'b01001000111010011001000011010010;
    #100 A = 32'b01101110000111110100110100000000;
    #100 A = 32'b01011100111011100110011110100101;
    #100 A = 32'b00010111001000100010010000101111;
    #100 A = 32'b00110000000111010000101100100001;
    #100 A = 32'b10011001111111111110000101101101;
    #100 A = 32'b00110111010101111100100011011001;
    #100 A = 32'b01110001100111110011001100011011;
    #100 A = 32'b00011100100000110001100100011000;
    #100 A = 32'b01011101100011010010111010100011;
    #100 A = 32'b00000111001000011010111011101100;
    #100 A = 32'b11110100001111100001000111000111;
    #100 A = 32'b00111111001010100010111010100001;
    #100 A = 32'b00001010100101010110101000101100;
    #100 A = 32'b00000001101110011011010011011101;
    #100 A = 32'b00011000010110111010111111111001;
    #100 A = 32'b01101110001011110001101110001000;
    #100 A = 32'b00000000100100001001101000111010;
    #100 A = 32'b00110010011101110111001110001001;
    #100 A = 32'b11000100001010100110101100101111;
    #100 A = 32'b10110000001001000010001001110111;
    #100 A = 32'b00010000110010111010100110011000;
    #100 A = 32'b01101101101111000111001000101010;
    #100 A = 32'b11110000111010110010110010010110;
    #100 A = 32'b01100101110001000101111101100000;
    #100 A = 32'b11101100101101011001011001110011;
    #100 A = 32'b10011001100100111001010010100000;
    #100 A = 32'b10111010101001100011110001011111;
    #100 A = 32'b10000010001011111110000100111001;
    #100 A = 32'b11101100100011100111000000101000;
    #100 A = 32'b01110010110110101000110011111010;
    #100 A = 32'b11101010110001110100100100100000;
    #100 A = 32'b10011000001111001001101110000001;
    #100 A = 32'b11100100001001100101010000110010;
    #100 A = 32'b10010100100000010111110111011100;
    #100 A = 32'b10101110010011011001110101110110;
    #100 A = 32'b00110001010010010100000100111011;
    #100 A = 32'b11000011100100001011010110001110;
    #100 A = 32'b10000111000111101001010011110100;
    #100 A = 32'b11011111010010111100110111000110;
    #100 A = 32'b11110011000111000101010101110001;
    #100 A = 32'b01011101001100100100000110011011;
    #100 A = 32'b00101101001110111101011100010110;
    #100 A = 32'b01110010100100001100011111101001;
    #100 A = 32'b11010100111001001111000011101000;
    #100 A = 32'b10011110010100001000011010111101;
    #100 A = 32'b01010011110000100010011010101011;
    #100 A = 32'b01011101001111000100111001011100;
    #100 A = 32'b01010001011101101001100001111011;
    #100 A = 32'b01100101000100000101101110010000;
    #100 A = 32'b10000000001010100011010111100110;
    #100 A = 32'b00010110111110011011001010111011;
    #100 A = 32'b10011010111101101001111000111101;
    #100 A = 32'b11110000010100101111011110011101;
    #100 A = 32'b01100011010111111001101111011101;
    #100 A = 32'b00010011101011011011111111001100;
    #100 A = 32'b11010001001100000000101011110111;
    #100 A = 32'b00100100000001001000010000111001;
    #100 A = 32'b10001100100100110001000010010111;
    #100 A = 32'b01000001000101011101101011000010;
    #100 A = 32'b11111001110000011101110011011101;
    #100 A = 32'b10110001011110010100011100111000;
    #100 A = 32'b11111100110100000111010100000010;
    #100 A = 32'b01000001010101010011111111111001;
    #100 A = 32'b10000101000100010010001101000110;
    #100 A = 32'b10010111100101010011111000011000;
    #100 A = 32'b11101010101000110110011000100111;
    #100 A = 32'b00111101000001110001101100001101;
    #100 A = 32'b11100100110111000111111010111100;
    #100 A = 32'b11000100010101111111001110000001;
    #100 A = 32'b10110111000110110100010000111111;
    #100 A = 32'b11101100000100011011001010111001;
    #100 A = 32'b11000110010110110100010001110000;
    #100 A = 32'b00100011100001101010101010100101;
    #100 A = 32'b01010011111101110111000110111010;
    #100 A = 32'b00000100111011010000110000010000;
    #100 A = 32'b11011010000110111111000000110010;
    #100 A = 32'b00100010101000111100010001011001;
    #100 A = 32'b00010111111000010011111010011000;
    #100 A = 32'b01100101010011101100101001010001;
    #100 A = 32'b01011001101011101011110101000110;
    #100 A = 32'b01111011011111111011010110111101;
    #100 A = 32'b11101010001001011110100101111011;
    #100 A = 32'b10111000111111011101000101010001;
    #100 A = 32'b00000000100111111001100011000010;
    #100 A = 32'b11011000110101101011001101011001;
    #100 A = 32'b11111110001001011100100000000111;
    #100 A = 32'b11000011011010111101010010110000;
    #100 A = 32'b01110111111011111101100011011110;
    #100 A = 32'b00000010111001110001011111110001;
    #100 A = 32'b11001111010110000000100011010100;
    #100 A = 32'b01000010001111011000110100110011;
    #100 A = 32'b11110101101100100100100111110101;
    #100 A = 32'b10000010000100011100110001100111;
    #100 A = 32'b11000001010010100110000001100001;
  end

  initial
  begin
    B = 32'b10100011111100110111101011111000;
    #100 B = 32'b01101010101001110011100100011010;
    #100 B = 32'b00100110110111111100001101011110;
    #100 B = 32'b01101010110110110010101111011010;
    #100 B = 32'b11111101101101111111110100100000;
    #100 B = 32'b10110000110100111110011100010001;
    #100 B = 32'b11110010001011000111110111011111;
    #100 B = 32'b10101101011100110000100010100111;
    #100 B = 32'b11011010101110000100001001111000;
    #100 B = 32'b00001011001110111110011000110110;
    #100 B = 32'b11011011000010110001110010011010;
    #100 B = 32'b11010110011110111100000001110111;
    #100 B = 32'b00111010010000001110011101010011;
    #100 B = 32'b11110010100101000111010010011110;
    #100 B = 32'b00000101010010100111000001110111;
    #100 B = 32'b01011011000000000100010000111110;
    #100 B = 32'b01110010001111111001101000101100;
    #100 B = 32'b00001110000001101111010001100111;
    #100 B = 32'b10010001000100110101010001101011;
    #100 B = 32'b11100010110000001110101100010110;
    #100 B = 32'b01011010011011100100110110100010;
    #100 B = 32'b10100001001000111101111000101010;
    #100 B = 32'b10000011100100101000010111010001;
    #100 B = 32'b10001010110100100110110010100111;
    #100 B = 32'b00011101001111010110010111010111;
    #100 B = 32'b11010100010001000001011001010011;
    #100 B = 32'b10010001001001110111010111111110;
    #100 B = 32'b10101001000000011010001000110010;
    #100 B = 32'b11110001110000111111000110100000;
    #100 B = 32'b11101011101010100010000000111011;
    #100 B = 32'b01101001010100000110110111111111;
    #100 B = 32'b11001111111111100001010101011010;
    #100 B = 32'b01001010011000100101110000110001;
    #100 B = 32'b00110011011100101010110010000001;
    #100 B = 32'b01110011011001111110000001010101;
    #100 B = 32'b01011000010100110110110111001010;
    #100 B = 32'b00010001110111101110011001110001;
    #100 B = 32'b10000011000100011111000100110111;
    #100 B = 32'b11010000001101111110101000100101;
    #100 B = 32'b11110101011000100011010010101011;
    #100 B = 32'b11111001111100110001010000010000;
    #100 B = 32'b11110010000001101000100000000010;
    #100 B = 32'b00000100100101010000010111110100;
    #100 B = 32'b10000000010010100001010000101110;
    #100 B = 32'b10110111111001111010001000100000;
    #100 B = 32'b11111110101101011001001111101000;
    #100 B = 32'b10110000000100011001111011110110;
    #100 B = 32'b10011110001001111001010001011000;
    #100 B = 32'b11100001001011010000001010101101;
    #100 B = 32'b10000100001101010010011101110000;
    #100 B = 32'b01111010000110111100101010000111;
    #100 B = 32'b00100001011111000011111011110110;
    #100 B = 32'b11011001110111100011111110101100;
    #100 B = 32'b00111000111000110101101101011110;
    #100 B = 32'b00000110011101000001010010000100;
    #100 B = 32'b00001010001011011000101110111101;
    #100 B = 32'b01010000000011100001111101100001;
    #100 B = 32'b01111010110110110011011001000000;
    #100 B = 32'b00010010100100110101100110011011;
    #100 B = 32'b01100010011110101011011010010110;
    #100 B = 32'b01100001111110001001101101100111;
    #100 B = 32'b10100001110100101010101101101111;
    #100 B = 32'b01110001010001101101100001111111;
    #100 B = 32'b10000011000100001010111011111111;
    #100 B = 32'b01111111100011001100000010101111;
    #100 B = 32'b00010000110111010100010011101110;
    #100 B = 32'b10011001110101011111010110100110;
    #100 B = 32'b11101101100110100000000010000110;
    #100 B = 32'b11000011011011001100011100010010;
    #100 B = 32'b11111101010100011110101111111100;
    #100 B = 32'b01101010001000100000000000111010;
    #100 B = 32'b11101011001010110100001010111010;
    #100 B = 32'b00010100010010100101001000001111;
    #100 B = 32'b11011001010010001010100101001110;
    #100 B = 32'b11101000011001011011010111100110;
    #100 B = 32'b10001110111001101000111111100111;
    #100 B = 32'b11111000100011101111101111111101;
    #100 B = 32'b00100000011110100000111000000000;
    #100 B = 32'b00100010101111011000011011101011;
    #100 B = 32'b01000110111100001110001001011011;
    #100 B = 32'b10100111111101010011100011000010;
    #100 B = 32'b00000011110111001011010101111001;
    #100 B = 32'b11110011010001000001110001100101;
    #100 B = 32'b10000000100000010001010101111100;
    #100 B = 32'b00101011110110111110110100000010;
    #100 B = 32'b11101101100101001101001011010010;
    #100 B = 32'b11110111000110000101001011010111;
    #100 B = 32'b01110111010000100000001111011111;
    #100 B = 32'b01100100100010100000011100011000;
    #100 B = 32'b11101100000001101111101111100000;
    #100 B = 32'b00110001101101011001000100111111;
    #100 B = 32'b10011011000110000001101110110101;
    #100 B = 32'b10110000110100001101101110011000;
    #100 B = 32'b01100101110000000000001101010111;
    #100 B = 32'b00101111011110101011001110000010;
    #100 B = 32'b10100000010111101011110100100001;
    #100 B = 32'b01100011101011010100110100111000;
    #100 B = 32'b01100000010010101010110101111111;
    #100 B = 32'b11101100001111000000010110001101;
    #100 B = 32'b11100110111000101100100110111010;
  end

endmodule
