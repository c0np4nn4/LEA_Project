module LEA_test_tb;

reg [127:0] Din;
wire [127:0] Dout;
reg [191:0] Rk;
wire [127:0] p3;

LEA_test
 U0 (
  .Din(Din),
  .Dout(Dout),
  .Rk(Rk),
  .p3(p3));

  initial
  begin
    Din = 128'b01001000000010010101110000010001011011000101011111011111010010111110011110011111001010011000010001110000110101001100000101001001;
    #100 Din = 128'b11000111101111000001101111011010010010001110100110010000110100100110111000011111010011010000000001011100111011100110011110100101;
    #100 Din = 128'b00010111001000100010010000101111001100000001110100001011001000011001100111111111111000010110110100110111010101111100100011011001;
    #100 Din = 128'b01110001100111110011001100011011000111001000001100011001000110000101110110001101001011101010001100000111001000011010111011101100;
    #100 Din = 128'b11110100001111100001000111000111001111110010101000101110101000010000101010010101011010100010110000000001101110011011010011011101;
    #100 Din = 128'b00011000010110111010111111111001011011100010111100011011100010000000000010010000100110100011101000110010011101110111001110001001;
    #100 Din = 128'b11000100001010100110101100101111101100000010010000100010011101110001000011001011101010011001100001101101101111000111001000101010;
    #100 Din = 128'b11110000111010110010110010010110011001011100010001011111011000001110110010110101100101100111001110011001100100111001010010100000;
    #100 Din = 128'b10111010101001100011110001011111100000100010111111100001001110011110110010001110011100000010100001110010110110101000110011111010;
    #100 Din = 128'b11101010110001110100100100100000100110000011110010011011100000011110010000100110010101000011001010010100100000010111110111011100;
    #100 Din = 128'b10101110010011011001110101110110001100010100100101000001001110111100001110010000101101011000111010000111000111101001010011110100;
    #100 Din = 128'b11011111010010111100110111000110111100110001110001010101011100010101110100110010010000011001101100101101001110111101011100010110;
    #100 Din = 128'b01110010100100001100011111101001110101001110010011110000111010001001111001010000100001101011110101010011110000100010011010101011;
    #100 Din = 128'b01011101001111000100111001011100010100010111011010011000011110110110010100010000010110111001000010000000001010100011010111100110;
    #100 Din = 128'b00010110111110011011001010111011100110101111011010011110001111011111000001010010111101111001110101100011010111111001101111011101;
    #100 Din = 128'b00010011101011011011111111001100110100010011000000001010111101110010010000000100100001000011100110001100100100110001000010010111;
    #100 Din = 128'b01000001000101011101101011000010111110011100000111011100110111011011000101111001010001110011100011111100110100000111010100000010;
    #100 Din = 128'b01000001010101010011111111111001100001010001000100100011010001101001011110010101001111100001100011101010101000110110011000100111;
    #100 Din = 128'b00111101000001110001101100001101111001001101110001111110101111001100010001010111111100111000000110110111000110110100010000111111;
    #100 Din = 128'b11101100000100011011001010111001110001100101101101000100011100000010001110000110101010101010010101010011111101110111000110111010;
    #100 Din = 128'b00000100111011010000110000010000110110100001101111110000001100100010001010100011110001000101100100010111111000010011111010011000;
    #100 Din = 128'b01100101010011101100101001010001010110011010111010111101010001100111101101111111101101011011110111101010001001011110100101111011;
    #100 Din = 128'b10111000111111011101000101010001000000001001111110011000110000101101100011010110101100110101100111111110001001011100100000000111;
    #100 Din = 128'b11000011011010111101010010110000011101111110111111011000110111100000001011100111000101111111000111001111010110000000100011010100;
    #100 Din = 128'b01000010001111011000110100110011111101011011001001001001111101011000001000010001110011000110011111000001010010100110000001100001;
    #100 Din = 128'b10100011111100110111101011111000011010101010011100111001000110100010011011011111110000110101111001101010110110110010101111011010;
    #100 Din = 128'b11111101101101111111110100100000101100001101001111100111000100011111001000101100011111011101111110101101011100110000100010100111;
    #100 Din = 128'b11011010101110000100001001111000000010110011101111100110001101101101101100001011000111001001101011010110011110111100000001110111;
    #100 Din = 128'b00111010010000001110011101010011111100101001010001110100100111100000010101001010011100000111011101011011000000000100010000111110;
    #100 Din = 128'b01110010001111111001101000101100000011100000011011110100011001111001000100010011010101000110101111100010110000001110101100010110;
    #100 Din = 128'b01011010011011100100110110100010101000010010001111011110001010101000001110010010100001011101000110001010110100100110110010100111;
    #100 Din = 128'b00011101001111010110010111010111110101000100010000010110010100111001000100100111011101011111111010101001000000011010001000110010;
    #100 Din = 128'b11110001110000111111000110100000111010111010101000100000001110110110100101010000011011011111111111001111111111100001010101011010;
    #100 Din = 128'b01001010011000100101110000110001001100110111001010101100100000010111001101100111111000000101010101011000010100110110110111001010;
    #100 Din = 128'b00010001110111101110011001110001100000110001000111110001001101111101000000110111111010100010010111110101011000100011010010101011;
    #100 Din = 128'b11111001111100110001010000010000111100100000011010001000000000100000010010010101000001011111010010000000010010100001010000101110;
    #100 Din = 128'b10110111111001111010001000100000111111101011010110010011111010001011000000010001100111101111011010011110001001111001010001011000;
    #100 Din = 128'b11100001001011010000001010101101100001000011010100100111011100000111101000011011110010101000011100100001011111000011111011110110;
    #100 Din = 128'b11011001110111100011111110101100001110001110001101011011010111100000011001110100000101001000010000001010001011011000101110111101;
    #100 Din = 128'b01010000000011100001111101100001011110101101101100110110010000000001001010010011010110011001101101100010011110101011011010010110;
    #100 Din = 128'b01100001111110001001101101100111101000011101001010101011011011110111000101000110110110000111111110000011000100001010111011111111;
    #100 Din = 128'b01111111100011001100000010101111000100001101110101000100111011101001100111010101111101011010011011101101100110100000000010000110;
    #100 Din = 128'b11000011011011001100011100010010111111010101000111101011111111000110101000100010000000000011101011101011001010110100001010111010;
    #100 Din = 128'b00010100010010100101001000001111110110010100100010101001010011101110100001100101101101011110011010001110111001101000111111100111;
    #100 Din = 128'b11111000100011101111101111111101001000000111101000001110000000000010001010111101100001101110101101000110111100001110001001011011;
    #100 Din = 128'b10100111111101010011100011000010000000111101110010110101011110011111001101000100000111000110010110000000100000010001010101111100;
    #100 Din = 128'b00101011110110111110110100000010111011011001010011010010110100101111011100011000010100101101011101110111010000100000001111011111;
    #100 Din = 128'b01100100100010100000011100011000111011000000011011111011111000000011000110110101100100010011111110011011000110000001101110110101;
    #100 Din = 128'b10110000110100001101101110011000011001011100000000000011010101110010111101111010101100111000001010100000010111101011110100100001;
    #100 Din = 128'b01100011101011010100110100111000011000000100101010101101011111111110110000111100000001011000110111100110111000101100100110111010;
    #100 Din = 128'b01011011111101110101110111110011000001111111100110000000010011010011111000100011111001001011101000011111111000100110010100001010;
    #100 Din = 128'b01001011111000010100001101111011001001001010001011000111010000011001001101101001101100001101001101011111010000100001011100111011;
    #100 Din = 128'b10011101101100001001101111011001111000101011000011111111000000111010000100101010000100101110010011110000001001011001100011110101;
    #100 Din = 128'b00010001011100000000001100010000011111010010001010100001011110011000110100111000111001001000100100111001110011101110100010110111;
    #100 Din = 128'b11001110100110000001001001110010110011101001110111100101000010001001010001100000110010001100101000010111011010001011010101110011;
    #100 Din = 128'b00011000000011100110010110010000010001001111010011101011110101010001010100110001110010010101111110001001011110110100111010001010;
    #100 Din = 128'b01011010011001110010000011111000001110000001100101000100101010001111011111001101010000000011001101100000001101001101101001100110;
    #100 Din = 128'b01001111010100101101110010110011000010011010000010010010000110001011100000101100011010111010100110101001001111100110111100101011;
    #100 Din = 128'b11010101010010000111001100001011101111101001000111101000011111010011111011000011111101010100110101111001100010111001011011011110;
    #100 Din = 128'b10110110010110110100110001110011110001101001001000010010001101100100111110111000111100001000000010101001011111001001001111100011;
    #100 Din = 128'b11001100010110101100101001000010000011010110010001111110110000010101000011101001010100000101010000101011111001101111001001111101;
    #100 Din = 128'b01100110110110000111001111100001111111010010000011100001010001101110011100111011010000110010100010001011101101111000001000100000;
    #100 Din = 128'b10100110001001011011000100000011111100011000101001000100010110100110100001011110111100011110010001010010110010111110001001100001;
    #100 Din = 128'b01110100100100111110011100011111110110101111011111011000011011111000100100100010001100011000110101110000101001101110111001101001;
    #100 Din = 128'b11011010111010101100010110110000111110100001001111111100100100101001011110111101110101000100100001101010001001001100111101000010;
    #100 Din = 128'b00010010000011110111010000000011001110010100111101101101101100111110101010011111010011110010011100100001100100100100111001110110;
    #100 Din = 128'b11111111111010110001111000110100010001001011010000001010111010001100010010100100111111010110100010001100101101111001011010000001;
    #100 Din = 128'b10111101110111011101001101011001111000100011111010010101001101011101111010101001011111010001010001010101011010110010101011111001;
    #100 Din = 128'b11000000011000000010010101001110000111010111000101111100010111100110100001011111000111000011100010001001011000001100011011000000;
    #100 Din = 128'b10100100110101100100110110001001011010001100000101100101000111101100011111001010110010101010011100110110111010010010100100101111;
    #100 Din = 128'b00100010001111000110100110110110011110010100110111110000111110111010111101011110111110111010110000001001110101000110100101000010;
    #100 Din = 128'b11010010101001110101010010011110001001010100000110010011010000001111100001000101110100110110111011111110111011011110011110111011;
    #100 Din = 128'b01000000100111010001111110010101110011111010110100011000001100011110100001110110110100011011010000000001001111111001010011010010;
    #100 Din = 128'b11100110110100000011000010010111111001001111011011010100101011100000001110101011110000010010001101000011110101110101101001000101;
    #100 Din = 128'b00100000001111110000000111011110001010111000111110110000000010111110010101111100100111001001100101010101010011101111110111000000;
    #100 Din = 128'b10011010100110010101101001100011010011100000110111111000011101000011010110001100101011110011111110010111111001011110011110001000;
    #100 Din = 128'b11000111010100000111001111001001001111000100110010100101011011100101111110110010111001110110111000110101011010111110001110110111;
    #100 Din = 128'b10101010011011001010100100100101001110100011110011110011010000111010110001110010010101010100010100101011010011000110001000001101;
    #100 Din = 128'b10010010000100000000001010010100111010010000001111101001000000111011010001111001101100100010001011001100101000111011000100010110;
    #100 Din = 128'b00010110111111000101011110111011100110010010100101110010101100001000111100100010111101111000011010001011001001010000101110001001;
    #100 Din = 128'b11011101001110101110011101110010100111001111011111001000011111001111011000010111001101101000111001101011100100011111001110101010;
    #100 Din = 128'b00010010110111111101001101111001000100011111001101111000001010101101111101101100100111100100011010100100001000010101001100001111;
    #100 Din = 128'b11110011100110010011101011101000000101001000000101100000001000011100101111000110111011101101110010011001000101111011010110000011;
    #100 Din = 128'b11100111010111011101010000000101100101101000110011111101000010001000001010011001110100101110101010010010010010111001101001100010;
    #100 Din = 128'b00000010101010011000101011001011110010111010000010101001110111011100001000101010110011010110000110110110011111101101101001001111;
    #100 Din = 128'b10111100001100100001000000011111101011010001001001000100101101000100101101010001101011010010101100100011101001111010110011010111;
    #100 Din = 128'b10100111100111000110010001111111000111100010100011110111001111101101110000111010001100101100100010101101000011000110110010101011;
    #100 Din = 128'b11111010000000101010110011100110101110000000001000010010100111100000010100111100111101011111010001000111000100100000111010010011;
    #100 Din = 128'b00011111100111101011000100001001001111110000000011111000110001001010010001000011101010100001010000011111110101111111010110110010;
    #100 Din = 128'b11111010101101001011101001111001000010110011000101000111011011111101111000101010111011010110001101111110011001111010100111101100;
    #100 Din = 128'b11011100000111111000000011001100000110000111000011101111111000001101000100010011010100111110110100000000011110101111011110000111;
    #100 Din = 128'b00001000011111000000000010100101101100000101011011011001011010011000110010001001011011000101001101011011100100011101110100001001;
    #100 Din = 128'b01010001101110000100000001011001100010011101011010000010101010100000000101000110100000110011100000010010001101011011011010111010;
    #100 Din = 128'b11001000100101001111011011010001101001111011110001110001000111110110001110101000110111101100001111001010111110101110100100100010;
    #100 Din = 128'b11100100011100100010100111100111010100010000100010111011111110000110000111111111101001010000001000010000110001110001000011110000;
    #100 Din = 128'b11001111010100001010010001110100110100100011000111001001010111100100111101110010100000101101100000111001110011101111111010000110;
    #100 Din = 128'b01110101101011000100100011110001010010011111000000100011110001110011011101011110001001010100111110011010011111111001010110011010;
    #100 Din = 128'b10101000100100111100111010001001101000100001100000001001100101011010100101000010111100100111011100001001001011010011100010100000;
    #100 Din = 128'b11010100001110111011100111001100110110001011010111100101001000100101100110011000111111000010110001100100100001110001101011001001;
    #100 Din = 128'b11101001100011011110000011100100000000101000010000100110010011010011101110001111010010110001110101011100101111101010110110101111;
  end

  initial
  begin
    Rk = 192'b001101111100110110110000110110000100000011101010001110010010000111011111110100100101000010011110011001011100011011010011111100111100000001001000010110000101111111100001111111111011010011010110;
    #100 Rk = 192'b011111110110010101100010000001000110011111110100101010100100110100011001101111000000001110011000111000111010011010100111011111111001101010100110000100100000010011111010011110001010000011101001;
    #100 Rk = 192'b000010111010110101001001101011010101000000110010011110110100110010100010000101001010100010011110011110000010110000101101010000011110101100100010000001000010011101100000011001001000001101110101;
    #100 Rk = 192'b110110000100101100101101110101101101111010001101101110110110111001111010101111111000010111110011110010000011000101110111111111100000111001101101110101101001101101001111011111101000010110000001;
    #100 Rk = 192'b011110010011110101100101111111010101111100101110100010101011100001100101011100011010110101111001110001000111001000010100101010100100011100100000100101100001110001110100010101010010011011101100;
    #100 Rk = 192'b100110110101111101100110100011110010100010010001001101010000000010110000011011100110101101010111001101001101000000110101001001101110001010010001111111000010000101100000011111011001001111010001;
    #100 Rk = 192'b111111100010110010010011000100100001110010001000010100110110110110000010000001101010001000011111010011111001100011110011010011000001101011011111111000010101001001011111010011010000100111000010;
    #100 Rk = 192'b100100111001000101100101011111001110011000001010000001111110000101010001111111110111000111010011011110010011111000011111100101111100001111001110110011100010011001101101101000001101010001001101;
    #100 Rk = 192'b100110011101001101110110000110011111000011010010000110110101111001101110100110010111010000011110000000100000101110011101101011110000010000001010001111101101011011000001001110001001101000000100;
    #100 Rk = 192'b100101001010101110110001001111111011010111010100110110111011010100100101010011001101101100100000100100001001000000111011110000000100101110110100010110011101101111111101001010111011100000010101;
    #100 Rk = 192'b111111000100001110111001111110110101011010101001010100000000000000001010001011011110010100100000000100001100100000001000111111101001101001111001000001010011111010011100110100110011001000010000;
    #100 Rk = 192'b101110011010000001011111111001101010101101011000110110110010110110110110011011001101111110101110101001111010000010000100101011100011101111100010110101001001100101010011010011100001000100011111;
    #100 Rk = 192'b000101011000100010001001001100100110011011111010111011000000010101001001100111100110101100001011011101100011010100111001011111001110000011000111000001110011011100101110011101011001011110100000;
    #100 Rk = 192'b001011101000011010010010010001110001100011010111001100000110101101001010111100010111100011110000110011100001110111111001110011111101110110111010000100100101000110101000000001110111101110100001;
    #100 Rk = 192'b001110111111101110111000100101000000000001001010110001100001011100010110111000001110010100110001001100010011111101100011010100010100010111001001111101101011110110010000010001000100010000100010;
    #100 Rk = 192'b101010111100110011101110000101111111000010111010101011111010000011101000011011011010000110011010010010010011001000000101110000000010110011000110100101010011000100001100010111001001101000111100;
    #100 Rk = 192'b000001100101010101001010011001101100011010001010000000001001000100100011110010011010101011111010100111100110011110110110110111100111010101001001100010110010110111001001101011101011000001111010;
    #100 Rk = 192'b001000000010110010111111101110101110110110011011111011110110111100001010111010011111100001100000101110010011101001001001001100101011111000011011011011000001001101000111010101101010001101010110;
    #100 Rk = 192'b011000101100011100010000100111011010100000110010111100100111110110101000010000111101101110111110000001011101111111010110111000010110011111100000001110111010010111000100110010011101011111001110;
    #100 Rk = 192'b110001100101000000011011111110100010011110000001011101110111110001011111110100011000101010000111110111010100000111111101100110100000011101010011111111001110110001110011110101000001001100001011;
    #100 Rk = 192'b011010010101000001000100010101101001111000101011001001111101001010110000001101111100111101010101111111100011011000100111110110101000111111000111101011110010100100101010010001011000111100101010;
    #100 Rk = 192'b000101000001111110001111100101101101110110011000101010110101100111110100111100010010000101010000101101000001001010110100111001001111111110111010110001101100010101010101001111010001000011110010;
    #100 Rk = 192'b111101111100111010101001110011100001000111010011100001001010101100111110011010001000000011001101110001011001110001010001100010100101111000011000100011000111111001010111011001001001100010110111;
    #100 Rk = 192'b110101111001010100011011110110101100110000111101101000110101001010101101001001010011001011101011101111001101100011100000011000010110101011111010001011110010111111001001100101000011001000010010;
    #100 Rk = 192'b000111001101001111011100110000111011100011001111101100100000111001110000010011111110000111000010101001001100001000111101101101111000010110010100111110011011100010111010010101001101001010100101;
    #100 Rk = 192'b001000000000011011000000100011100100110010000001111100110011111101001110011000000110111100010001101110001100011110101111001110111111011000101010100010000110111011001001000000110101101110100100;
    #100 Rk = 192'b111100111101111111100011010100000110011010110100001111001010001011110000110011001100101111100110100100001100110001110000010100110001000100111110000010100001011001100000110010101111010001101010;
    #100 Rk = 192'b111000000011110011000101100100000010010111110010000011001100000000111011001100111111111000011000000011101101011011000100101011110100100000111101110001010000011101010000111101011010001010010111;
    #100 Rk = 192'b000101011000001011101000101111111001011111101111110111110011110110100101111101001111100000101101111011011100111011100100100000011111010011101001101001100110100101101101100001100011011101011111;
    #100 Rk = 192'b011010010011001010000110001001010100000100101000111010001111100110000000010010010001010000000110001101000111000011111101101000001000001010011010000001010110100010000101111100001110111101100000;
    #100 Rk = 192'b101010001100011000011110100101110000101000011111011011110111100011011101110011101001101101000101010100011010010111111100001011000111011111110001110011101000111101001110011101110110111011110011;
    #100 Rk = 192'b110110100010110001101001000011110100001111010010100101110000110101100001110111110001001101011111100111111010100100011001111101110100011100000110001001011000001001110111111100010001100010010010;
    #100 Rk = 192'b001110000100010011000010001101111011110000111101110101000111000010010010011001001111000011011110010101010001111110100111001010110110011000110110111110000100110100110111011011001000001011110101;
    #100 Rk = 192'b110100010110101100011110000000101011101110000001101000110001001001001001101100000001001000110111100111101111000001001111101111100011101000001100000111111010010010001001111110010011110101000000;
    #100 Rk = 192'b101100110100101111111000011000111000011000000010110100100110111100101010101101011001001010110000011001001000001001110111100100111010100110101100110100000000011011111101011110111110111010010111;
    #100 Rk = 192'b111110110010101001001101010100010010001111010000101011010010001011101000000110011100110010101010011010111000100101000110110110000111011101010110111101111101011001010110110000000001000110111110;
    #100 Rk = 192'b011000001010010100101010110100111010010101100001001101010000011011111000001010010100110001001001000110110110011101100110110110010110000001000110010100001110001000110111100001110010100011000001;
    #100 Rk = 192'b100001111101110111101100010010111100011110110100111010100000011010001101100010111010100110000100001000111011010001110101101111100000101011000000110100100011101000011000100001001101101111110101;
    #100 Rk = 192'b111110100100110100110010000011011010001100001010000100001000011100000100000000001111101011111001101111110010110110000000110101010100110000001000001110011011001010011011000101001001101001101110;
    #100 Rk = 192'b010111110001101000100110011001111011000011111110010101101101111010100011011000010110001111111110010101001100000100010111101001101000111110001111010110000000111001010010111010101010001000110001;
    #100 Rk = 192'b100001110011011000000010110110011100101010010110001100010110011110001010100110111101100011000001001010111111011000011111101000011011110111110100111001000011101101011000100010111011110000101001;
    #100 Rk = 192'b100011001010001001011100101100000101101101010100000100000110110000000111001101010000011011010010010111010001101001000101010111000100111000000011110011110110000010101100100000100001101110010101;
    #100 Rk = 192'b100010000010001011000001110000000000110101011001100010011010110011010010101011110111001101011011001000110111100110001100000011110011111011110000010111000111101000010000100011001000010110110110;
    #100 Rk = 192'b000111011001101101110111011101110000000001111111011110011010111111011011011001100101110110101100010101111111101001000001011011010010110001111010111000100101000101011001111011111101110110000001;
    #100 Rk = 192'b011010001010110011000010001011000100000110111010001010001101011001001000110100111110111000000110110101010110100101011010011011001011010000000000100111110100000011111001000111010001100011011101;
    #100 Rk = 192'b000010110110010100101000111010111101111011000011001111011111110110100010010100000110011101001101100001010011011110000110011100110001000001111000111001000111100101000100111111000000110000111111;
    #100 Rk = 192'b101011000110100011011001010000001111001100011110010000110001000110000000001010001100111011000101101011010011000101010010001110001011001011111110101100001001100101101100010101101010110010100111;
    #100 Rk = 192'b110010101101101110010110100000110110110100000011100001100001101010001010011000101100000001101000101110010011110001011010001110001001001001000101001100101101000101110001100000011011111101101011;
    #100 Rk = 192'b110101111110000110111011100000100100110101011011100100011100011001001000011111111010111000111011111011011101100000000101101011000110101000001111100100000001111110010100000000101001000010110111;
    #100 Rk = 192'b011011100100010100010110001010110100001111010010011010111100001010110111111100000011001110111110100001010101110100011110011010010011111001110001101001110111011000100101010110100111010101110110;
    #100 Rk = 192'b100011010101101000101001010011010111001111101001000011100100000110000001010010110001111100111000000010111100001100010111000000100111100000010111101101011000110110110100110010011001101110110011;
    #100 Rk = 192'b001011010011000000101010110110010111000011101011100000111000110100000010011001111111101101000110000001101100001000101001111110000111011100111011100110011100000000001000101100010000111000111000;
    #100 Rk = 192'b101011010000101010010011001001000100010111000110110110000011011000101100100000101110000001001001001100101100011000110010101101000001101010100100011110111000010111100111000010010000000011010011;
    #100 Rk = 192'b010010110001111011111100011111001010010010001101111011111110111110110000101110001100100001100100001011000110010111001011011000001001000010000100110111111111110111101000100100001101101101111101;
    #100 Rk = 192'b100100101100111010100000110011011101101101110011110101110001110110101100111001010010011110101101011111111110110100111011010101101100101101011011010111111101110001000111101110101011001001101111;
    #100 Rk = 192'b101010111001011111011010011100001001100101001001110101001101110111010000101000110001101010000110011011000010100110111000010001011011011010111010100101011010011000001001010100001100110101001111;
    #100 Rk = 192'b010101101101000111100101110001111010000100011010010010000011110000011100110011110001111001000000001101110101100110011111100000010110001100110000100000110011010011011100010111011111000111001101;
    #100 Rk = 192'b000111011110110001001000100110001100110000101000101000001001111100010001000001110010100010111100010100001110100010101001110100111010110100011110110100010100000001010011010101111011011101001000;
    #100 Rk = 192'b110110000110011000100111010000011001001011001111010100000101100110000100101010010100100100011110111000011100101100110100000010110000101010001000001110010101101011111100101010110101001100111010;
    #100 Rk = 192'b011000100100111111111110100100001111101010111011111001111111111101010011111001000110011001001001110100111000100111010100001110100110101110110111001101010111101000101100101000000101100010111100;
    #100 Rk = 192'b000001011111111010111010100000101110110101010110011111101000010010111100001111100000100101001001011100111111111011000010110001100011101101010010001110010101101101100111101101100000110001100011;
    #100 Rk = 192'b001011011111100111001011000111000101000111000000111011111100001000110000101101001111011110010111010100111000101011110001010100100110000010110001101100100111111111010110001001010100101001100011;
    #100 Rk = 192'b010111100101110101110100010000010111111111001010111110011000101001001101100101110110111101001111010111010101100001000111110011110001110011000001100010100101111000111111101101111110111101010100;
    #100 Rk = 192'b100010010011100100011100101001010001011000010110000001000001010001011011100101001101110010101001000111101010100100010100000000111111100110000100011011111101011010010010100010011010001011111000;
    #100 Rk = 192'b100100011001100001100011011011100101101111000001111110100111110001110101110110011010000100010100111101001000110000010000111110100001011001010001010100111000100111000111011100001110110110101100;
    #100 Rk = 192'b100011100010000110111100100001010100011100111111010001010101101100100011110100011100100111101111110010011101010000010101001010100010111001100110100111011111001011011101100010011110110110100011;
    #100 Rk = 192'b001101111110110101011001101001001011001000001010011010100000110001111111111111101001101110101111111100111101101111011000110110100011011110101101101001100100011011100000000100001100101010110000;
    #100 Rk = 192'b001111101000000100011100010011111000101001000011111011101100101101101111110111100001011101100101100000010001111111101010110011111011001010011101011001101010010010011010110100011011010000100000;
    #100 Rk = 192'b110110010100010000010110110110101111001111010011011001011011000101001101000110001000010010001111010000111100011111110100001010101110100110011100100000110101001010111111111000011001011011100111;
    #100 Rk = 192'b010001110111001111110000100101011111010001101111011111010001110110111011100111101001101001110011111110010000010110100110111010111010110110111000101000011011001011010111100110111000101010011001;
    #100 Rk = 192'b010110110010011011010000001101010011110001101001111110110100000111010110110010001001011000100101000011001000001010100000000010011000010011110011001000101110010111001110110100111110110011100010;
    #100 Rk = 192'b100001011001100101111110001010000011111110100110101110100100110010101100110111010111010101000011100010010011101000011010100001000101001111100011001001111001111001010000111011111101011011000010;
    #100 Rk = 192'b111000000110101011111011101010100101011001010001110000000100000110111101100100000110011110000101010000101010110110011100011011111010101001101100101011110000011111101000110000001111000000110000;
    #100 Rk = 192'b110001011101101011101111000100100010101001010010000011011100010010000100000110101010101110111110011000100011111100110000001010011001010100011110101100011001111100101101000110100011110111110010;
    #100 Rk = 192'b000111111011110010100110101111101101110001100101000000010001011110110111011000001001000011110100110100011101100111000011001111100011101000101111101101000101000001111001101111100101101010100010;
    #100 Rk = 192'b011111110110100100001100110000010111011111100011001000010000100100100110100101001111011100110011001010101001101001101000110010111011101000010011110000011001111010101110000011011010010110101111;
    #100 Rk = 192'b001100111000111111110000010111001010011100011000001100010001000001110000101111110101100111100011110110101011010111111110110000011110100101100111000010000010001101011101001011101101111111111110;
    #100 Rk = 192'b101101110010110100100001010010010101110111001000011011001101100110011001100110100011010111101111000001101100000001010011010100000110011011011000111111011101011110001010100101100010100110010100;
    #100 Rk = 192'b100100010010111000000011001111010101001101001010011111010111001101000010111100001011011010001111001110100100110111110110111101110001000101011011000011100000100001101100100110010110100011000110;
    #100 Rk = 192'b100101010100011100010110011001110011001100011111110001001000110010110011101100010011011101000000010100010000011000010011110010100001101000000110100011010101010110001110101001110100101010111110;
    #100 Rk = 192'b011011000110001111001110100111000000010100101010100111011100110000011011010000000110100101110101010111001010000001111010100111010000010111110011101110111101010100010111010111011100101010011001;
    #100 Rk = 192'b000100111000111000100011000011111100000000100100000001000011001001011110001000011101010010101000011110100100010010110110101010010100100100011011111100011101000101101000101110100010101111011100;
    #100 Rk = 192'b011010010100010001110111100110001011011111110101000011001110110010110110000011011111000110011000010001100111110000111111101000100101010000001100111010110100011101111110101000001010101110000011;
    #100 Rk = 192'b100110100111010101011111011101001100101111000110110001111100001010011100010110000011001010001010011110010111010000100100001000011001001011010001000011111001001101111010011010110111000010100110;
    #100 Rk = 192'b100110101000001111110101001100100111101011101110100111010100111010111011001110010001000000010110011000011010001000000110111001110011010000011001000100010111101100001000110011010110011010100010;
    #100 Rk = 192'b101010011111000000000001001100010001100011011000111110001101101011111101101001000010000010100000110111011101101111101110101110110110011100111101001011001110101111111101111100111101100010011000;
    #100 Rk = 192'b101011111101001100010000001011111110010100001101000010000001100111110000010111010000101011010001010011100011101001011100100101011011001111011001001110110000100111000011101000101001000001110100;
    #100 Rk = 192'b100100000001100010100101100110111101010101111001001101101111110100101010111101111001110100011110100000011110110010001100101100000110000011110101001101111100111010011100101000110110100100111001;
    #100 Rk = 192'b000000001001110000100000111101101011000101110100110011000100110100101001101010000110010110010010110011100110110001011111011111101111101000010100110100111000110001001100101101010110010001010110;
    #100 Rk = 192'b001001101001011110111000110100011000101101001100101000100001101101011110110101001111111111011111000110101111111001110000111101110001010101001101011010101001010101000010001000111000000110011101;
    #100 Rk = 192'b101001001000110011011101111110100101011001100001101001110100010110110011111000101010011000111101101000111000001100010111100010111110010101101001010010111111011011111110101010001111110101111000;
    #100 Rk = 192'b100100000111001010100010000001000001101101010100001000110100001000010110001011110100011001011010100001111100000001110101010011111110011110111111110110001110110011111001101011101100000111110000;
    #100 Rk = 192'b000100010010000101001100101110000010100000110101000000011011001000001010011100010101001010011001100010101100011001100110010000010111101001001011001010100101001010100111111101001010101000101010;
    #100 Rk = 192'b100000111010111100001111011101100110111000100111011100111000010110000100010000001110001100111111100010111011011101100111111010100011101000010110100111100101000010011111100000111111110101001011;
    #100 Rk = 192'b001111011111010111111111000101011010001010000000000110111001110000011011001111101111001010100101010001011111101001101101100010001100100101001100110000011011100111011111111000100011111101110001;
    #100 Rk = 192'b001111101100000010101101011011001100001000101010101011110111101010111001011101110111011011010001110000011011100001100000001001011010000100101001111010101111001110111100000000001100100000011110;
    #100 Rk = 192'b111011100010011100100010001111110011001000010011101101100011011101001101011000011001011110111101111101100101001011101101011010101100000100001011101010101001111010110110110101001100000101011101;
    #100 Rk = 192'b110000111011101100011001010100110100111000100100000001010110101010100100011100101001000010010001011000011101101011101101011001110111010001000000001100001011100110110100000011010111000110010100;
    #100 Rk = 192'b000111010011101111101101100110101100101111110101101010011111010001011000000110101001100001101011100111000010010011001011111010010100000000000011111000101000111100000110000000001001101110001010;
    #100 Rk = 192'b111100111110010100011100001010111000001110101001010110000011111100010110011110001101111010000010110001011010001010000111010100110001010000000111101101001001011101110001110011010111001111110110;
  end

endmodule
