module LEA_Encrypt_tb;

reg [127:0] Din;
wire [127:0] Dout;
reg [191:0] RoundKey;

LEA_Encrypt
 U0 (
  .Din(Din),
  .Dout(Dout),
  .RoundKey(RoundKey));

  initial
  begin
    Din = 128'b11000011001100110101111010010111100011101101001001001110100010000100110011010011001101001010100111000001111101010011000011101110;
    #100 Din = 128'b11010111101111010100000100000011010111000101101011100011110100010101100000110011001100011000111110101000001111100010110110101110;
    #100 Din = 128'b11101101111010000100110011000010111101100111000000100100010011111111101111110011101000010111110010000010110100001000010110110000;
    #100 Din = 128'b11110011001111100011001011011011001010000001011110100010101110111011110101001010001011100000110001011110010000111111110000011101;
    #100 Din = 128'b00100111100010010100111101110010110101100101100110101011101010110100110101111000100101011001110000111000000110111010101001111100;
    #100 Din = 128'b10011100101011010110111100100000101011010010011001100100001100011000001111110101000010110001101111001000001011101011111001010011;
    #100 Din = 128'b00001110011010101111010110001100110100100010010111111000000110100000011111010011010101001110000101001100000101110111010010110101;
    #100 Din = 128'b00010010101110011100010111110000010000110100110100111000101000101011010010001111110101000110111010011001100100110001001101110011;
    #100 Din = 128'b00001111101100101011001000110101111110001011000110010010100100100111001111100011010100001111000101001111010111101110100101111101;
    #100 Din = 128'b11100011100010001010000011100101100001101001001010001111101011111001010100100011001101111101011100111010010000011011011011000110;
    #100 Din = 128'b00110011001001101010011100001101100010011110011111111110101010101010110001110000000111111001011101011111111001100100001100100010;
    #100 Din = 128'b00100111001010111110000001100000001011001111100010010001010001000010110101110011100011101001111111010101110111000100110101011100;
    #100 Din = 128'b11011011010101110011001011001101001111000010000011001010001010010000010111110111000010000111110100001111111101000011100001001110;
    #100 Din = 128'b01001110111011011001110000110110011010001010010010011111101101010101110101010010110111101010101001100001000010001111001010101100;
    #100 Din = 128'b10111111001111101110100101011100010110100010000011100100011101111010011101101001110110101010010010110110010111100100001010000001;
    #100 Din = 128'b01011010011000110001111011011001100110110001001111011111001101101100010011100000100000010110000011010011101000110000111111001000;
    #100 Din = 128'b01101110111111100100001001100010001011100001000111100101001100001010011010001100111010101101110110101110100010000100111100010101;
    #100 Din = 128'b11100011001111001100010110101000001010110011110000001111111000111100000110011101001101101111101110111010111111001010101101101000;
    #100 Din = 128'b01100011000110110110100100010001011110100100001111101111000000100101111110010111000100010101101000111011010010011010101100100000;
    #100 Din = 128'b01011011100011100000011000111001010001010001011010010110101011011000010101000000011101101111010111001000001100001101000001110010;
    #100 Din = 128'b11111111010011000111111001001000010110101011001001000001111101111111110010010000001000010011100001101001100100101011000011011011;
    #100 Din = 128'b01110100100110101100110100110010011010000110101000111010001000100000011001000001101011000010110001110110110011100110100101010110;
    #100 Din = 128'b11011001100100011111101010001110000110001110100110101010111011100000000010010101000110010001110101110110010111110111100010110101;
    #100 Din = 128'b01110101110110001111100100001011000100001000011111011100000011101101110010101101101000000111110001010010001010111010101111100010;
    #100 Din = 128'b01010110101111101001110111011111100011100011100111001011010100110010000000010000011111101010011000101011111001010001111100101111;
    #100 Din = 128'b10110101000011110110011111010010101011101010110010010010000001111010111101111010000000011000000000000110000111111001110110010011;
    #100 Din = 128'b01000011000110001010110100011000110000010011110001100111100100000100100010010111101011010010000101010100110011101000011001101001;
    #100 Din = 128'b11110000010110101100111110110010001000001101000001110001001111000101000100001011100110010010101101011010010100111110000100110100;
    #100 Din = 128'b01010111001111110110110001010101110111110101000010011010011001110100101010101110011100011101011110111100111101001110010100101101;
    #100 Din = 128'b11111010001101111010110110011010000010111101011110110000110000111101111001010111100011100011100000000000001111010100100111101000;
    #100 Din = 128'b10111010010000010100101101010000010000001010011110100101001110010001000101010010011011111010111100000111000100101000111001011011;
    #100 Din = 128'b01101110001001100000011100010011110011001100000011010101101100000010001100111010110001100101001010110010101110110110001001100110;
    #100 Din = 128'b10110011000100001011011011110110101101111101101100101001010111110111101101011111100110001111101100100111101110111010010100010110;
    #100 Din = 128'b10100101010100111100100110110001010110110100110100110000001101100101000111000010101011000001101011100110111100101101011110011001;
    #100 Din = 128'b01000111011010111101100101001010001111010111001110000011010000000110111000010111100100000000101000000101100111010100001110110010;
    #100 Din = 128'b11010000001011010110001000101100000110100101010110101001110001000101111000101011000100010010001010111111001010111100100100010110;
    #100 Din = 128'b00110001101001001000111000001110110100000100001101010111110101101100010001011011001001111010111110100001001001010011010001100101;
    #100 Din = 128'b00111100110101011010001010000010110001010111101010100110001101000010111101011001111001000100010001111011011100110110010111110000;
    #100 Din = 128'b11111000001100100100010111011000101101010010010111001001111000101011001110001100000000011101001010011011101001111011111111111110;
    #100 Din = 128'b10100010010001100011010011011010101011011011111111100101101101101101110001010100100000010010100100001001000011111110001010111001;
    #100 Din = 128'b01100000100101001111010011011101001000001101100011110001010000110101111000100110011100100100100001011100001000001001101010110010;
    #100 Din = 128'b10011111011100010110011010011101111111101011100000101101111101001001101001011101111010001101100101010011101001010110010111110110;
    #100 Din = 128'b00001111011111111001100000011101001101101100001011011001110010110011101011001010011110101000110100101010110000101111010010111010;
    #100 Din = 128'b00011001011100010110110001011101111001000100101011111100011001011010100110101001101001110011000101001110111100001111000110111001;
    #100 Din = 128'b01011100101101010100111100011001001001110011000001111110011110101011100011001011111101100110000101111001110001110100111001000100;
    #100 Din = 128'b11111001011111101100101101110101111101011010000111101110111010111101000011001011001001111010110110111100110010000000100100011100;
    #100 Din = 128'b11000011111000100101010111110011101101111100001000110100011010110011010110101111100000011101101101000110101000111101110001101001;
    #100 Din = 128'b01100101001111111100111111011000101010001110001001110101000101101110011111100110110110111101111011100101000010101111011001110011;
    #100 Din = 128'b10010101110000010000100101101001111111111101111010110111010101101010101000100110001001001010001011100001010011111010100111111010;
    #100 Din = 128'b00011100001011000001110000101011011001000001000011011100110111110110001000111001101101011100010110011111111010010100010000111101;
    #100 Din = 128'b01100100000111010100110010010000010011001100101011101001111101110110001001110010011100001100011010111010001100010111101011001011;
    #100 Din = 128'b10110101000011001101010011101111100110101100010111001010101100010000000101110101011011010001100011110110000110000001110110011000;
    #100 Din = 128'b10001110000111111010101010010101101111000010010001000111111100111001111100011110010001011011101010011100111001000101011111100000;
    #100 Din = 128'b11110011010101110100001111111111101010010111010010001100000100011100110011001111001111000011100011001111001000101010001011000101;
    #100 Din = 128'b11000110000000100111111001101011000100000111110110011010100101111111110000010110110110000111100111101011101100101000010110011010;
    #100 Din = 128'b11110001110011111111101011010011111001010010111000111111001001101111011111110100111000000000010001110101000000111100101110101001;
    #100 Din = 128'b11111111001010110100010100000000001000101100010011111010011010011100001101000001011001100100010010110011000101010101011011010011;
    #100 Din = 128'b00111010110100101111001101011110101111011110111100110100011110100100000010000000000111110010010011001110111011110001101011110010;
    #100 Din = 128'b00010000000011010010001001110011010100100000001101110000010100100011010011110001100000011111110011100000001101111001010110100100;
    #100 Din = 128'b00100100110011111001011110010101001001001111001000001100010111111101011101111101101011011011111011101111100000110100100001101010;
    #100 Din = 128'b10101100100111110010011010010111101001011000001001101101011100000101011110111101101110000101110000110101000000101000110100000000;
    #100 Din = 128'b10100111011010010110010110001010010111110111111001010100100011101001011101000000000010011001011001100001011010010100001101011011;
    #100 Din = 128'b10011111000110000111001101111110011000011001000101000010111111100000100000010110011000001001010001001111010101111010001111000111;
    #100 Din = 128'b10100011001111001100000000010110001111100011110100011111101011111110001000111111000110100000010001111101010110101110011110101000;
    #100 Din = 128'b01110000111111100111000110111010011110111110010101101100000101101000001001101001010000101110011100000010111111000000000001001111;
    #100 Din = 128'b10110100000000111000010001110110001010000001111011100111011011011011111011111100001110000001100010001010000101110011010111101111;
    #100 Din = 128'b00010010000010010111000011111010100110100100010011010110111110000001100000110111011010111111000101101100010101000010001001010000;
    #100 Din = 128'b01010010011101011111000010010001101001000001001010110001101100010011101011111010011111110101100001110110111101111010010110001110;
    #100 Din = 128'b10111010010110110100111000001101110111000000111101100001111001011100101100010011010111010010001010000100101100011010010101111101;
    #100 Din = 128'b11110100000001001110100001111111011001001110000100000001010110111011001100101001100101100010001010010101100011111000001001000001;
    #100 Din = 128'b10101111111110001111000111011110000110100110010101011111001010000100011011101011011000011001010101001001000001101011001011111000;
    #100 Din = 128'b01111000101010001101110101100101001111001011101000001111110111010000011110000001100100111011011011100101110001110011010101100001;
    #100 Din = 128'b11001001101001000011101101001011011000111011101001010110000110101111011100000111111100011010110111000011010110100100011110100111;
    #100 Din = 128'b11000001001110101011011110110011101000110010110111011101101110101001011110111000010000000111111011110000111001011111111110100011;
    #100 Din = 128'b00100000011110100011010101001110010110101101010110011000011011011010001010110101011110100010101111110111111001111111000000111011;
    #100 Din = 128'b00111011011101000011000001101101110011100010110011010001001001110100010100000110000001111001111101010110100100011110111010011100;
    #100 Din = 128'b10010001101100011000110101111001110110101110101110011110001111101010110001001101010110100110101111011010110011011011011000101011;
    #100 Din = 128'b11001010101100000011110101010111001011001011111100101100101101110011000111000100111101111010110000010011110111000011110110110101;
    #100 Din = 128'b00110111010100011111100111010111011111101010101011000101111101100010101100101111111110110111101111111010011100011001010100010101;
    #100 Din = 128'b01000010101010100001000000101010000011100101001111101110011010101000111001110010100100011000001111101101111001101110110100011111;
    #100 Din = 128'b00011110010100110101100010010111110100001101011100010000001111100111100110011100001110111110100100001010010100010001011001011000;
    #100 Din = 128'b00100100010100111000010110000110111001000001111110010101100001111011010010001000100000110110100111011101100011011111111000101010;
    #100 Din = 128'b11011011011111110110110001110010110000011110110100111100111111001010000110011000111010100000111101101010001101000101111100101010;
    #100 Din = 128'b11000100110010000001111100000101011011010001110111000100110011111001010000000110001100010000110001110111111101010100001110111001;
    #100 Din = 128'b11011101011101001111111011110100000001011100111100000000100001011011000000010111011011100001010101010000110111111101100010000011;
    #100 Din = 128'b00011011011000110011011100010100110001100010110101111111011010110011100100001011010100100111100111001100101010111111000101111111;
    #100 Din = 128'b01101111010111001111001101101010011100111101010110011010001101101011110011110101111011100001000111010000100000011011010111111010;
    #100 Din = 128'b01000000101001010000001011001101111111001011101100000001001010001100010010111011001010000001100010011000000111100100111001110011;
    #100 Din = 128'b11011001110000011000101110111101101010100010111100001010011101110100100011101100111101011110001011010100111010110101011001000001;
    #100 Din = 128'b00011000011001000001001100001001100110001100000110010101100011100001001110101101101100110000000111111001101100100111010011001100;
    #100 Din = 128'b11100010101101001011100001110000001100111100010010110000111011111111110100101010100101011111111010101111101100111010101000100010;
    #100 Din = 128'b01111111010101101001100010110110100000010100110010001111001011110100001011000111011110010110011100011110010010100000010100111110;
    #100 Din = 128'b00010100100110111100011010111100101101111111001110101100001101000011010001100101011010010111100111111110000100001100101011001101;
    #100 Din = 128'b11111100001110101100011110001010110011000011100011000100111100001000011010100011110000001001101000110101111001000100000110000010;
    #100 Din = 128'b01100111001100011100010011010111110011110001110110110000011100000101011000110100100011001011011000001001010000001011110010001000;
    #100 Din = 128'b00100000100101011111001101001101110110010101010000010010101101011101101010101101000110001100110110011000000000101110101101101101;
    #100 Din = 128'b10100001111010111011011111100101011010100000100001111101010010001100011101110111110011100010001110011010110111001111101110101011;
    #100 Din = 128'b00100101111000010101100001101011001010011011001010101101101111000000100111100000000100010110111101110010111011111011101111100110;
    #100 Din = 128'b11001001101000111111000000010100011000101010001101000111010100000010000110111110011001101010101110111010110111010001000010110000;
    #100 Din = 128'b11001000010101110001010101011000111000000011110001001010011011001110001100111110110101100100110001101010001010101110000111101001;
  end

  initial
  begin
    RoundKey = 192'b000101110000110000001001010011110100111011000000011001101111111100110110000101001010101010101110001010110011011010001011110101110111110111101100110111101011010111101000001100010010010110010010;
    #100 RoundKey = 192'b001110111000011111000101111110110101011001000010110000001001110010100100100111001100100000101110000100010111000101011110110011101100101000001110000110111001110010110010000010011101110011011001;
    #100 RoundKey = 192'b101110100110100101000111001101101110011010110111001111011111110001011110000110110110101110010111010010011010101010110000010100000010110101101001011000111101010100001010110001111111000101001111;
    #100 RoundKey = 192'b010010011011111000000010011000110100110000000010111010000101010001010000000101101000010100100110011010111011011101011010000011011010100011101011111011110101010000101110001001000001110111111101;
    #100 RoundKey = 192'b000110010000010010101110001010101100001111001110011010111111101111001000011100010111000000011011011101011111101001101001101111011110101110000001110000101101011100110010001011000000100100110000;
    #100 RoundKey = 192'b101110010001000001010010000001001011101110100101110011100110110100000110011001010111010011110000111111101101010101001110011100010010111110110000000110000000001110101100010010011110011110010111;
    #100 RoundKey = 192'b010010110000111111100000001101000011010100001110001000011010111000101000001010111010101001011011001011111011100100101010001010010101011011101000010110011100010010101111111110101011000100001110;
    #100 RoundKey = 192'b100011111000111100001100011010100101001010011100001100100111100000001000110001011111010100110110000000001011111011001100011111111001100101110011100101100010100101011011011000111111110010000011;
    #100 RoundKey = 192'b101010011101011110111110100000000011000110101011111101100010110111010100001110101000000110011100011110011110001111101000010101111110010110100011011010011111111101011011100000010110000001011001;
    #100 RoundKey = 192'b100010000000010010100110011100011110110011101100001001000001111110101000100100001100110111011101111100100101001010001011101101101011000111010001111001110011111001111111111010011011010111101111;
    #100 RoundKey = 192'b011111100010001000101100011111101100010110111110001101110010100110101101000101111000110010001111111001001111010100111111001111011001100001111011110001111100101111011100010101011011011110111100;
    #100 RoundKey = 192'b111010111010110010101110101110111001100011110011111010110100110110011000000100111101000010110000001100110101010101011011101101011000011011111010001100010100100100000101011111110000011111010011;
    #100 RoundKey = 192'b000001000100010001001000111000111011001100100101100111111110100010000111100100000000101111011001100001010100100101011101110000101110101000001001111011010011100000101001010111100101101000101000;
    #100 RoundKey = 192'b010110010110110110011101100110001000001010010110101110110111101011010110101101001000011110000000001001111110111100101111011100011011111110110101100111111011110110011000001100010000101101001001;
    #100 RoundKey = 192'b011000101101110111111011101111111100101111110101100010011001001011000010010000101011101111111000000100101101001010001111100100111101000110000100100000111011010001011100011101010001010100011010;
    #100 RoundKey = 192'b101101010011001000010100001001110010001011110010000111011110100101101101011101010110110011111110110101001100011001000110001100110101000001001001011110001100010101010101010011111001000011001100;
    #100 RoundKey = 192'b110100000100101010001110010011001101111100001100011010110100110000000101000000111111111101100110010110110111001010001010001011001001110111010001101110111010001010101100001101011000110110001010;
    #100 RoundKey = 192'b111101111100101000011011010000100101000001011000111000110011010010101110110110100101100010011101111101111001010101010010111110010011111101010100110111100000111110110000001101010111111000101111;
    #100 RoundKey = 192'b010001010111010100010001001000000000010110011000101001011001011001101110000111011111010110000101011001000001001100011000001100100000101010111001010101010000000100001100111001000000110101111000;
    #100 RoundKey = 192'b010100101100110000100000000101110000011000110010011000101011011110011101110010001111001010111101111101010111100010001110111100100111111111001001100101100101111011111110101000101011011110110100;
    #100 RoundKey = 192'b010110001000111001001011010100001011101110100110000101111000100101101111100011000100101111101011111000100011110001101110110011101111001100110000011011110100100101111110000101111111110000110101;
    #100 RoundKey = 192'b111100100110101000001011011000101011011101000111010011110101011100001010101001101111010001110010001100101000111111011000101100000001010011111001101101010111101100110011011111001010011010101010;
    #100 RoundKey = 192'b000001101101100000101100010110010110010011000100000111111110111111100110111001111011000010101001011111000000101110000000011011110010010100100010010000111011110011001110011111011101111000110011;
    #100 RoundKey = 192'b100110101010010111101100111010111101111011011100101011011101011011110001001101110011100111110000111111111001001110100011100011110010001101110110010011010111010010011001111100110101110000011010;
    #100 RoundKey = 192'b010111010100011000011111110111001101110111001011000000100011101010011110001111101011001100110110001011010101010000110001010111000001011000000001111110001010111100100110010111001100001101110110;
    #100 RoundKey = 192'b000100010000000111001000101111001000110110011001100110011001100111100011000010010010111100011110110100111111100101010010111110110110110010101110010111001000110000100110010110011100100100000101;
    #100 RoundKey = 192'b110100000011110111100010100011111110110100111111000111001100010101100101000010100100110110010100000110110010100000101010111001000010101001110101010101001110110010110011110110001000101100001010;
    #100 RoundKey = 192'b101101000000101010011000000111011100001111110111100000110101110001010110011100000110100001110011010111101000111001100011000011011011001110110111011001101100010000100011001101001100100001011100;
    #100 RoundKey = 192'b100001011101100101001101101001010100110110110110010110101000011010000111010001011110001111010000110000100111110110100000101001100000011110101001010011100101000010100001101000110110111010110011;
    #100 RoundKey = 192'b111101010110010101010111010000110111011010001010111001111001101101110111001010011100101101000001001010001000000100011100011101001100101101001101011111110110011110001111111000110111000101011000;
    #100 RoundKey = 192'b001110011001110000001110111110111011111010101011110111010000000011110000111001001011110001011110010000100111110110001101000011100011011001010001011101101010101011010111010010001000011000000000;
    #100 RoundKey = 192'b000101000110100101001111010011111110010100110010011101100100101010101010111100000100001110100100101001011110000000110101010110110101011001010110010001001001001100010000100100000010110010010010;
    #100 RoundKey = 192'b101010000000110110101011110100100000100000100100001010111111100001110110110011011011000001110000001010100110110011110110100100010010010100111011111100000000001101010101001000000101010011001110;
    #100 RoundKey = 192'b010110011010000001110011101010101001011011111010100101111001000101110101011111101101000100011010101011000101010110101001111001011100011111010111110100001001010010000010100000010011100110001100;
    #100 RoundKey = 192'b011101000110111011011000001001011101000111101111110010101100011000001100101101010110000100110001111000100111111111010100010101001110000001110101010011000001000011110011111001111011000110001110;
    #100 RoundKey = 192'b110001101010100100111100100011011001101110000111000111110110001011101100011000110101101001010111111100101100111011000101001010100001101101011100100011111111010101011001111001111001011110010000;
    #100 RoundKey = 192'b101011010000100000110011111001101001110101001110011110001011100011110000010100000010010011000011010010011100110101110111110100001001001101111001011011000111010101001001001000110100010110110111;
    #100 RoundKey = 192'b111001011101111110111111010101001000010010011110000011110010101000010000111001101100111001111010010111110101011010110110001111000101111011111111001011101111111111000001010101100111001000001111;
    #100 RoundKey = 192'b000010101000011000001101010101101010001100101000011100000001011110000001110011001110011100101100001011101100000101010001110100111011100111000111110100101001010101111111000001011000100001010010;
    #100 RoundKey = 192'b010101001101100010101010110000001100001000111100011010000001110111100010110010001010111101000011111011101101011100010101000110100001111011111100010000001001001010101000111101100000011100001001;
    #100 RoundKey = 192'b110111111000001110000001101110011110100101011110101100101111011000100110101011100011000111111100001110001011010010100101101101111011101110011110101001011001111110111000011001101100000001100011;
    #100 RoundKey = 192'b111111101000000110011000000100000011101110100111110011100100001000101111100000000110000110000100111101110110110100011000110101000010000100010001111001111000010110100101101100110011010001011000;
    #100 RoundKey = 192'b000111011100011001010010001000010100011110011111001111101000010110111001101111110011011011010000100110110001001000011001100011111001101100001001110011100101110011000101011001011100100011010110;
    #100 RoundKey = 192'b011100010110001011110000110100010011011011110111001001001011011111111001110011000011010001001110110111001000101111000101010101101100001000111010110000110010111010100010001110100000011000000110;
    #100 RoundKey = 192'b010110000010010011111010011101110001100011001111001000100101010100100011111101100010001101101001110100101101010111011111011100111010000101001101001110111000100001011100111010100110011100000010;
    #100 RoundKey = 192'b110100100101010000100101101010101001011000100110001000010000111110000100101111110110001110101110111101000111001110111101100000110000110110000011010010000011011110000100011100101010111000001011;
    #100 RoundKey = 192'b001100111010100111111111001011100001001011101000110011011111010110011000101001100101101111011010001000011011100011010011010100011110011001001001101101111100101101110001000010111010000000011100;
    #100 RoundKey = 192'b011000000001000001101100010010101000100011111000101100110000001111010000111111101011011101101111001111010001100111101010110000101010010101000011000111100010101110101001000011010010011001000110;
    #100 RoundKey = 192'b011000010110000010100100000010010011100001010111011001110000100111010011011010110101110000111100010110010111110101111000110011100110101100111011100011000001010111111000011001111001001100100100;
    #100 RoundKey = 192'b101110110010110010000011100011010010001010011101110001111001100111101000011010111110100011100010001011001101101000010110110111100010011000001000000000001011010000011010001010010000001010010111;
    #100 RoundKey = 192'b011000000110000000000100011000011111000011001101010010001000101000000100100101000110010000111111110011000111001111101111101000111110000011000101111000111011001010001100111001011011110011011011;
    #100 RoundKey = 192'b011010101001101100011011110001010101101011110001100110100001101101101110000001000000111110110000000010010000101100000111100100101100100000010000101101011111011001111011100011001010011011010000;
    #100 RoundKey = 192'b001100001101111110100110100100001010100001100111011110011101111111100100010010101011111101000010100011100111011111111000000110101100010011000001010110001110101101101000011111101110000011001100;
    #100 RoundKey = 192'b010010111101001111100011110000101001111000010101010010010111001111010000111001101101010001110100011101000000001110110010011011010100101111110010010000000011101101100110000000101011001001100111;
    #100 RoundKey = 192'b010110100110001110100001000100111000100111101111010111100001000010011110101000010100111000101110111000101001011101111101000111000101011001000001101111001110011000110101000110100000010001000011;
    #100 RoundKey = 192'b110101001000000111011101011100001010001001110100011110010010100001111010111101001001011111110101010100001011100110001101001010101000010111011110111101001001010110100101100100001010100100100011;
    #100 RoundKey = 192'b110111000011111000111000000000110100000000001001011010001001010011101101110010011111000011100110111101111110101101100110010101111010111000110010000001001101010101010101101011000111101101001110;
    #100 RoundKey = 192'b001100110100011010101000000111000000110000111110110100100100100100101000010001101111001100101001110001111110100010110001101000010101000111111110100010001000110101111000010011011101101010010111;
    #100 RoundKey = 192'b110101000110000010111100101100100101001010011001111001110101000101001010001000111000001101001000111001001011001111110001101110010111000000011001111111011011000010001110111110110100110111110110;
    #100 RoundKey = 192'b000000101010000100001110111101010111100001000100100001100100111001011000000100011101010000001010010011000000000110111000100111010100001011011011110101000110100111001001000011001001111010111101;
    #100 RoundKey = 192'b000001100010111100110110111110111100001111001110110001100110110100000011100000011001110011000111001111101110111111001100100011111011111110111111111111100000110111110010001011100110011111001000;
    #100 RoundKey = 192'b001101100111111111001101111010101110101011011011001110100100111011100000010001110011111101101100101011101100011001011010101100100100100100010011010001010011110110011000011111010111111110110111;
    #100 RoundKey = 192'b101000111101001110100010000000000100001000101100100101001001000110001000000000010001001101011100110110111101111001111010001011011110001110000011000011101110110011010000110001111011011001111001;
    #100 RoundKey = 192'b011110101000100010010000111000100100001101010110000111000100101110010100101010101101010000101101001001010011010011111110011010101000000010011100110001011101011011101011100011110000101000111001;
    #100 RoundKey = 192'b110110010011111100000010111110000100110110100100010000100000101110101100110000110100100010011001101110111000111100111000011110100000101101000101111101001000101111111000110011101111111110111110;
    #100 RoundKey = 192'b110000100100000100101010110100010011100010010011111110001110100111101100100001000011010111101001001110110011111010011100110101100110011111101000110010101010101010011110001110110001101001011101;
    #100 RoundKey = 192'b110111100110101101111011001110100111010100110000100100101110010000010100000111100011011100001101001010001100000101001011011111101101010000000100011000111011010100111111110000010110000001010011;
    #100 RoundKey = 192'b011111000111111101010100001111000101000110110100101010110011011101001001110000111011111011111001110111101010011000100011001101101001110001010000001010100001010100010100011010011000001001001001;
    #100 RoundKey = 192'b100001101110010111000110011010001110001100011110011011010010100000111001000100101101010101100111100110110010010100010111101011110101111001111111001001111000100111011100010110110110000001011001;
    #100 RoundKey = 192'b011011000000010111110001010111000010110110111100111111001111001101100101110010001110011001001100111001010000110010001010110001110100010011100101111000001000011000101111001011000000000000110010;
    #100 RoundKey = 192'b100110011110000110100000101010100011001111001000110011011100100110011001100011001101100010110011000001001011010001010011110010001001101100110010000000001011111111100001100010011010101111110000;
    #100 RoundKey = 192'b101110001101110011011101111101000010100001100010101000100110101010010011000101010001001110011001111001011110010011001010001010010010110010010101011110101101001100101100001110100101010000011111;
    #100 RoundKey = 192'b001100011010111110101111010101010000000111010101101010000010111001010101111110101011101100010111100100001110111001011100010100111000110100010011000110001000110000100110110111011000101000110111;
    #100 RoundKey = 192'b110010000000000000111010100000011011000001111001001001100101110000011110001101000001000101111011101001000101111111000101110111011110110101010011001110001011001000000001000010110000110100000010;
    #100 RoundKey = 192'b011001001011111100001010100011110111100100011111101101000110101010000010010111100000011101101011011101100001000111100111101110001001111000110100010111100001010110010100010101000011111001100110;
    #100 RoundKey = 192'b011001101000101001101010110110000001010111100000101011111010110111111011110111110011100100110101011011110001011001111001110010011011111011010111000100101011101000011010100001101001100100101010;
    #100 RoundKey = 192'b000010101001110100001001101100101011110001111110110011000110001000101001111000100010100011010101111110001010001100101001111101011100001001010010100000100010010010101000101110000110000010101101;
    #100 RoundKey = 192'b001010011011010001111000010100001000011001010000011010110110001101111010100011111011111100110111011101100010110110000011000100111011011111110100101011001111110001001001001110000110001110011001;
    #100 RoundKey = 192'b000111011100110000000011001010111000100101111110100101010011011011111000011001011111101110100100011000100111101000110011110010100110100111100110110101111000010100010010101001111110110010010111;
    #100 RoundKey = 192'b001000101011001011010100010001011010001001001100000001100000101000110010110000100011001000111110001111101101101010111100111000011100001110010000111110010000110010011000110101100011011111101011;
    #100 RoundKey = 192'b100011100000100110100111100001101011000010010101100101000010101101101001000000101010001000101100110011101100011101111010110000100001001111111111111000101101001011100110010110100111101000110111;
    #100 RoundKey = 192'b000010000110111110010100001101000000011010110000000000101100111100010101100000000001100001100101101001001110001001111001011010110000010001110101111111001011101001110100011110110110110100000001;
    #100 RoundKey = 192'b100000010011111001011101100110001011111000010010110000100100111010110000010000100000111111000001000101000000001011001011111101001100010110101101111001001000011001100111110000101101000101000100;
    #100 RoundKey = 192'b101100101110110000110001111000001000001011010111111011010110111010100000101110000010101100010000100101010110111010001100000111010110010110010100101010011010101111101110111001111110111011101000;
    #100 RoundKey = 192'b001000011010100000110001110011011111001110101000100111000101100000001011000000110000011100110000011011000111001001110111010100001101010000110001001110010011100011011000110110101001100011100110;
    #100 RoundKey = 192'b100100001111100000110011010110110110101111000110011101000100011101101000011100001111010011000011011001111110111001110010100000011110110101111001010010111000110101010000101100011100011111010011;
    #100 RoundKey = 192'b000011010111010101111000110100000010110110100111110100100001110110101000101000010110010001000110100010100001111001000010110011010111000111111011101001101010011011101111110101110000010010101111;
    #100 RoundKey = 192'b000110100011111001101110011111001000110000101110111111001111011011001000001100010101111101110000001101101000010101101010010101110001000100101000001110110110000110000011101111000100000110010100;
    #100 RoundKey = 192'b110110110010100110000010101100100100000001100001110000100100101111011011010101010011111101001000100011011011110100111001100110110100000001110011000101010100000001000100001011010011010011001000;
    #100 RoundKey = 192'b111110101110111100001100010110110001100100111100111101101000111110001111010011011111100010000101110101011101100000001101011110111000001110011110100110111001110001000010101000110100100111010001;
    #100 RoundKey = 192'b011110100000111100101100010110010001100110000110010001100101100010101100101110100011111101001011100010110011010010011101000010110111101011000101010110101011110111010100110001110100101101010010;
    #100 RoundKey = 192'b010001111100100101111011010110011110000010110010100011110110110110010011000111101011000000110001010000111000010000000001111100000001100011111010010110101100100111100001100111010001010111111001;
    #100 RoundKey = 192'b001110101000011010111011010000100111000000000000010001101001110110100000110111010110100111101010110011110101001100110101110101111011010011100100001001110010101000101111010111000001000100101100;
    #100 RoundKey = 192'b011011110111011000001000100010010010101001111111111000000000011001111000100111111001000111111011100100010100110101100101101001010111100010100101111000100010100101111110110001100101111010101100;
    #100 RoundKey = 192'b110101101110110001111101010000011010100010010011111011001011110011010100000010101101101100010000000011001000010000100101100011011011100111011111000110011110111101011011101100000110100010001011;
    #100 RoundKey = 192'b011101000000011110111001100010111010010010111100001001000100101100001000100110001011111110101000110000001110110010011001100101110111001011100110010101011100011111011001101110001101011110100101;
    #100 RoundKey = 192'b100000001000011010101100101001110001000001000111010100011110011101100100100011110101101110011101000101011110000100010001111111111101110110110100000000110100110101000010111100101100010010111111;
    #100 RoundKey = 192'b000100011111101001001010000110110000111010001110000111110011111111101110110001101100110000011111100100010001111111001001011001100001101000010100010000010001011011100100111101110101011101110101;
    #100 RoundKey = 192'b001001010111010110101000000011001100010101011100001000000001010101101101001000011101100001011001011101001101010101100100100000010111111010110001010111101000001110111000111101010001100010001000;
    #100 RoundKey = 192'b100101000110000001011000101010000111100101111100110001101001101011101011111101000011100101000101100011001000001110010110110110111001010011010110110100001110100100000001101101110101000101101100;
  end

endmodule
