module LEA_BlockXOR_tb;

reg [31:0] Block;
wire [31:0] Result;
reg [31:0] RoundKey;

LEA_BlockXOR
 U0 (
  .Block(Block),
  .Result(Result),
  .RoundKey(RoundKey));

  initial
  begin
    Block = 32'b01011111111101010110100000001010;
    #100 Block = 32'b00100011001110010101001011010011;
    #100 Block = 32'b01110100010011000010010101001110;
    #100 Block = 32'b11001010000001110010001100100001;
    #100 Block = 32'b00011010001111011101110111100110;
    #100 Block = 32'b01010000011110100000011001101110;
    #100 Block = 32'b10101011110001100100100110011110;
    #100 Block = 32'b00101110110110111110000011001001;
    #100 Block = 32'b01111111001111000110010011111010;
    #100 Block = 32'b11101011001000101101011100101110;
    #100 Block = 32'b01000100001000101110011111110011;
    #100 Block = 32'b01001011001001110100101101110011;
    #100 Block = 32'b10000001001101110111100110010001;
    #100 Block = 32'b01100110111111100001000001010001;
    #100 Block = 32'b11001011111101110100110010101101;
    #100 Block = 32'b01101111000100001100000010101010;
    #100 Block = 32'b00110010000110110110101010110100;
    #100 Block = 32'b01101111001111100110111010111110;
    #100 Block = 32'b00001111001101111010000001000001;
    #100 Block = 32'b00110011000101100110011110010001;
    #100 Block = 32'b10110001010001110011111110111010;
    #100 Block = 32'b01010011111001100011101001100101;
    #100 Block = 32'b01001000111001010101000001010010;
    #100 Block = 32'b01111011011001001011100000011100;
    #100 Block = 32'b10011101100110110010011011111011;
    #100 Block = 32'b00001011101010000011001001110111;
    #100 Block = 32'b01100100011101111010001100010000;
    #100 Block = 32'b10001100011101011011000110111001;
    #100 Block = 32'b01100100100100011101111111111010;
    #100 Block = 32'b10001010101110000100110111110110;
    #100 Block = 32'b00111111101100000000111011001010;
    #100 Block = 32'b01111100010011110010101011100001;
    #100 Block = 32'b10111111011001100110110010110010;
    #100 Block = 32'b10000000001111101001011001111001;
    #100 Block = 32'b01111010110011101011111111111110;
    #100 Block = 32'b11100010100110101000010000001110;
    #100 Block = 32'b00001010010110101110000001000111;
    #100 Block = 32'b00100001100100000101001001100000;
    #100 Block = 32'b00100110011001110111101000100001;
    #100 Block = 32'b00001100001011001110001000010101;
    #100 Block = 32'b00101100111000000100101010110101;
    #100 Block = 32'b11101110101001101100010001011110;
    #100 Block = 32'b10111111000100000010001010010100;
    #100 Block = 32'b00110111110001001000111000010001;
    #100 Block = 32'b00001100110010101100111000000010;
    #100 Block = 32'b10001001110100101011111111010110;
    #100 Block = 32'b01000110110111110110110110111001;
    #100 Block = 32'b10110001101011101110100101110011;
    #100 Block = 32'b01011010101000001011110011010100;
    #100 Block = 32'b00101011111110011011111101010001;
    #100 Block = 32'b11010100101110111111000101011011;
    #100 Block = 32'b01110111001011011011110110000101;
    #100 Block = 32'b01001111001011110111111110100100;
    #100 Block = 32'b11111010101001010100101001010001;
    #100 Block = 32'b00110101000101100001101010111111;
    #100 Block = 32'b10110000110101110111100100110011;
    #100 Block = 32'b01000011000101000110000011000101;
    #100 Block = 32'b11110000111001100111010010111110;
    #100 Block = 32'b01010110010101110001010100001100;
    #100 Block = 32'b10011111111000100001000000110110;
    #100 Block = 32'b00001101100011101000101001010011;
    #100 Block = 32'b00000011110110011111101110110001;
    #100 Block = 32'b10011101011111000010110111011001;
    #100 Block = 32'b11000010000011000101110000101100;
    #100 Block = 32'b00110001111010100100110101011110;
    #100 Block = 32'b00111101111011111000100111001101;
    #100 Block = 32'b00010111101100000101011110101101;
    #100 Block = 32'b10011101110000111000010000110011;
    #100 Block = 32'b11010001100011100010001100100110;
    #100 Block = 32'b11000010000011010101011110100110;
    #100 Block = 32'b01101011101011000110110101001101;
    #100 Block = 32'b10000010000000111010101001010111;
    #100 Block = 32'b00111001111000101010011110100111;
    #100 Block = 32'b00100001111110111010011110110001;
    #100 Block = 32'b00000010111100010010001010111101;
    #100 Block = 32'b11010000100100101010000100011111;
    #100 Block = 32'b01111100100100011011001011011001;
    #100 Block = 32'b00001011111001111001101011010100;
    #100 Block = 32'b11011111111100101111001100100101;
    #100 Block = 32'b11111011010010101001100101100010;
    #100 Block = 32'b10000101000011100100011111001111;
    #100 Block = 32'b10110101010000111111111110000011;
    #100 Block = 32'b10001011101111110001001111101011;
    #100 Block = 32'b11001101101100101110110001001110;
    #100 Block = 32'b11010101110100001101000011100010;
    #100 Block = 32'b00101011011111011000100001101010;
    #100 Block = 32'b01110101101000101011100011101101;
    #100 Block = 32'b10111011001111111010001000111000;
    #100 Block = 32'b10100000010110100011110111110100;
    #100 Block = 32'b10111111101011011010101100101100;
    #100 Block = 32'b10110110000110000101101000010101;
    #100 Block = 32'b10010001101010001101011001011010;
    #100 Block = 32'b00100111101000000000011100100101;
    #100 Block = 32'b00010000110110100010011110110000;
    #100 Block = 32'b10000011101011111010001111000101;
    #100 Block = 32'b00110010101101101010011101111011;
    #100 Block = 32'b01010101101010010110011010011010;
    #100 Block = 32'b01001110000001001110001001111100;
    #100 Block = 32'b10110100101010100110110000011010;
    #100 Block = 32'b10101000100110100101000000010101;
  end

  initial
  begin
    RoundKey = 32'b11101100010110000001010110101111;
    #100 RoundKey = 32'b10000010011101001110100110000001;
    #100 RoundKey = 32'b11010111010011101010001101001001;
    #100 RoundKey = 32'b11010000001110000010010010100111;
    #100 RoundKey = 32'b01010010101111111101010011101111;
    #100 RoundKey = 32'b10001011010101000010101010001011;
    #100 RoundKey = 32'b01101110101011101000100100101001;
    #100 RoundKey = 32'b01100011100010010000100110011000;
    #100 RoundKey = 32'b10101000110001110100000111110100;
    #100 RoundKey = 32'b11110010100010010000111101011111;
    #100 RoundKey = 32'b11110101101100011011001100010100;
    #100 RoundKey = 32'b10000011011011001011011000111111;
    #100 RoundKey = 32'b00100000101101111011001100101101;
    #100 RoundKey = 32'b01110111010111011101001001110000;
    #100 RoundKey = 32'b11011100000111110000001110011011;
    #100 RoundKey = 32'b11101111110111010110101001100111;
    #100 RoundKey = 32'b01010101000111101000100110110011;
    #100 RoundKey = 32'b00011110000111111111100001110010;
    #100 RoundKey = 32'b11101111111100010000000110011001;
    #100 RoundKey = 32'b00101011100011000100111010001000;
    #100 RoundKey = 32'b00100110110100111100010110111000;
    #100 RoundKey = 32'b00101001101111100000011011001111;
    #100 RoundKey = 32'b01100100110001001100010111100010;
    #100 RoundKey = 32'b10111000110001101101000000010000;
    #100 RoundKey = 32'b11001101100101110011101111110000;
    #100 RoundKey = 32'b01000010111110100010100111010001;
    #100 RoundKey = 32'b10111110010110010111101000111101;
    #100 RoundKey = 32'b11100100101111011101110110010010;
    #100 RoundKey = 32'b11100100100001010111010010100000;
    #100 RoundKey = 32'b00100101111101001011111011100010;
    #100 RoundKey = 32'b01101000001101000100011000000001;
    #100 RoundKey = 32'b00111111011100111011010111101001;
    #100 RoundKey = 32'b01001111110111010011000001010001;
    #100 RoundKey = 32'b11100111100111101010101001110110;
    #100 RoundKey = 32'b00100001010010001011100110001101;
    #100 RoundKey = 32'b01010101110000110000100100001100;
    #100 RoundKey = 32'b11001001011101110010101100100000;
    #100 RoundKey = 32'b10101110101001011001101011100000;
    #100 RoundKey = 32'b01110001110011001100100111111100;
    #100 RoundKey = 32'b10100001010111001100111010010001;
    #100 RoundKey = 32'b10100011010011110001101000110000;
    #100 RoundKey = 32'b00101101100011110111001101001101;
    #100 RoundKey = 32'b10100111111010000110100101100111;
    #100 RoundKey = 32'b11100100111110000101101010000101;
    #100 RoundKey = 32'b00100010001100010111011100111010;
    #100 RoundKey = 32'b11110011100111010011010010101101;
    #100 RoundKey = 32'b10110111101101110011000101101111;
    #100 RoundKey = 32'b10011101111100100111101011101101;
    #100 RoundKey = 32'b00010111001100001101011111011001;
    #100 RoundKey = 32'b10101111110110000000110101000111;
    #100 RoundKey = 32'b11101111000000010101011110010010;
    #100 RoundKey = 32'b01010001110110001101110101000010;
    #100 RoundKey = 32'b10010001000101011100011000011010;
    #100 RoundKey = 32'b00001000001011100110100011010011;
    #100 RoundKey = 32'b10111110101111001111001101111010;
    #100 RoundKey = 32'b01001011000100010001101010111110;
    #100 RoundKey = 32'b00111110011010101010010101110101;
    #100 RoundKey = 32'b10110111100100101100110011011000;
    #100 RoundKey = 32'b11000101010100000101011001010101;
    #100 RoundKey = 32'b01101001010101110100010100011010;
    #100 RoundKey = 32'b10000001110000011101111111111111;
    #100 RoundKey = 32'b11111000010101011000110001111101;
    #100 RoundKey = 32'b10101100011100100100101011010011;
    #100 RoundKey = 32'b01101010010110111110110111001001;
    #100 RoundKey = 32'b01101000101000110000001100011111;
    #100 RoundKey = 32'b00111001101010001001110001101001;
    #100 RoundKey = 32'b00011010100011100000000101111100;
    #100 RoundKey = 32'b01101010010000011100100000001101;
    #100 RoundKey = 32'b10110001011011101100111101000110;
    #100 RoundKey = 32'b00111010011010011100010011110000;
    #100 RoundKey = 32'b11001101100100010000110101001101;
    #100 RoundKey = 32'b01011011100111100111101011000001;
    #100 RoundKey = 32'b10100111001110000000101110000001;
    #100 RoundKey = 32'b10110111000111010010010111110111;
    #100 RoundKey = 32'b10101001110101010100101110011101;
    #100 RoundKey = 32'b10010101001101111001110110010001;
    #100 RoundKey = 32'b10100101110111011000111110001011;
    #100 RoundKey = 32'b10010100110110111001100110101101;
    #100 RoundKey = 32'b10000101001010001101110100011100;
    #100 RoundKey = 32'b11000011011010011011100101100111;
    #100 RoundKey = 32'b11111111000111100000000110100110;
    #100 RoundKey = 32'b01101001111110111000011101100101;
    #100 RoundKey = 32'b10111010010100001000011010001110;
    #100 RoundKey = 32'b00101111100111110110110011010010;
    #100 RoundKey = 32'b01011100000011110001101011100010;
    #100 RoundKey = 32'b10100100000001100010111100111111;
    #100 RoundKey = 32'b00011011010010100101110011101010;
    #100 RoundKey = 32'b01100011010010011000110000000100;
    #100 RoundKey = 32'b10110100111110000101101000110111;
    #100 RoundKey = 32'b11001010000110111001000110001100;
    #100 RoundKey = 32'b01110101110010101111111100000100;
    #100 RoundKey = 32'b11001110011000000110001000110011;
    #100 RoundKey = 32'b00100000010001111100000111011101;
    #100 RoundKey = 32'b01010000101011110101101010111111;
    #100 RoundKey = 32'b01100011110100101010010001011011;
    #100 RoundKey = 32'b10100101001010101101000100110000;
    #100 RoundKey = 32'b00111001101000101101100110111101;
    #100 RoundKey = 32'b10011111100100001110100110010011;
    #100 RoundKey = 32'b11101111110010001000110110011111;
    #100 RoundKey = 32'b11101101110001111111101100110101;
  end

endmodule
